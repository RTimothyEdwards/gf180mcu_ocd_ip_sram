magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect -133 -66 160 595
<< polysilicon >>
rect -14 529 41 562
rect -14 -34 41 0
use pmos_5p04310591302060_512x8m81  pmos_5p04310591302060_512x8m81_0
timestamp 1763476864
transform 1 0 -14 0 1 0
box -174 -86 230 615
<< end >>
