magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< error_s >>
rect 4781 2303 4792 2306
rect 4837 1941 4848 2303
<< nwell >>
rect 5024 6624 5936 7070
rect 4666 5394 8559 5744
rect 4659 5194 8559 5394
rect 4659 4844 4666 5194
rect 4713 4080 8559 5194
<< pmos >>
rect 5231 6723 5287 6935
rect 5367 6723 5423 6935
rect 5544 6723 5600 6935
rect 5673 6723 5729 6935
<< pdiff >>
rect 5119 6920 5231 6935
rect 5119 6748 5143 6920
rect 5189 6748 5231 6920
rect 5119 6723 5231 6748
rect 5287 6723 5367 6935
rect 5423 6920 5544 6935
rect 5423 6748 5457 6920
rect 5503 6748 5544 6920
rect 5423 6723 5544 6748
rect 5600 6723 5673 6935
rect 5729 6920 5840 6935
rect 5729 6748 5770 6920
rect 5817 6748 5840 6920
rect 5729 6723 5840 6748
<< pdiffc >>
rect 5143 6748 5189 6920
rect 5457 6748 5503 6920
rect 5770 6748 5817 6920
<< psubdiff >>
rect 5727 7588 8460 7622
rect 5727 7541 5793 7588
rect 8385 7541 8460 7588
rect 5727 7506 8460 7541
<< psubdiffcont >>
rect 5793 7541 8385 7588
<< polysilicon >>
rect 5203 7111 5259 7127
rect 5564 7126 5623 7332
rect 5231 6935 5287 7111
rect 5367 7081 5623 7126
rect 5367 7066 5600 7081
rect 5367 6935 5423 7066
rect 5544 6935 5600 7066
rect 5673 7014 5816 7072
rect 5673 7007 5751 7014
rect 5673 6935 5729 7007
rect 6327 6998 6383 7126
rect 6246 6944 6462 6998
rect 6246 6935 6302 6944
rect 6406 6935 6462 6944
rect 5231 6672 5287 6723
rect 5367 6672 5423 6723
rect 5544 6672 5600 6723
rect 5673 6672 5729 6723
rect 6246 6617 6461 6690
<< metal1 >>
rect 4635 7588 8460 7616
rect 4635 7541 5793 7588
rect 8385 7541 8460 7588
rect 4635 7513 8460 7541
rect 5126 7173 5207 7513
rect 5282 7106 5364 7387
rect 5439 7173 5520 7513
rect 6241 7107 6323 7292
rect 6398 7221 6479 7511
rect 5282 7023 5520 7106
rect 4936 6920 5209 6945
rect 4936 6748 5143 6920
rect 5189 6748 5209 6920
rect 4936 6728 5209 6748
rect 5439 6920 5520 7023
rect 6241 7014 7205 7107
rect 5439 6748 5457 6920
rect 5503 6748 5520 6920
rect 5439 6673 5520 6748
rect 5753 6920 6240 6938
rect 5753 6748 5770 6920
rect 5817 6748 6240 6920
rect 5753 6738 6240 6748
rect 6316 6743 6397 7014
rect 6472 6738 6756 6938
rect 5753 6729 5834 6738
rect 5439 6589 6438 6673
rect 5948 6470 6042 6589
rect 5388 4009 5479 4391
<< metal2 >>
rect 503 7586 594 7679
rect 751 7586 841 7679
rect 1647 7586 1737 7679
rect 1900 7586 1991 7679
rect 2789 7586 2879 7679
rect 3036 7586 3127 7679
rect 3951 7586 4041 7679
rect 4177 7586 4267 7679
rect 5578 7357 5668 7451
rect 5189 7249 5435 7337
rect 4984 7014 5846 7108
rect 5016 6649 5134 6873
rect 5928 6647 6046 6871
rect 6639 6642 6757 6866
rect 5948 4542 6038 6481
rect 5588 4448 6038 4542
rect 5588 2853 5679 4448
rect 5748 3585 5837 4391
rect 6572 3868 6662 4391
rect 6932 3444 7022 4391
rect 7115 3187 7205 7113
rect 7756 3727 7846 4391
rect 8115 3303 8206 4229
rect 5786 1648 5877 1742
rect 6970 1648 7060 1742
rect 8154 1648 8244 1742
<< metal3 >>
rect 4753 6803 8515 7384
rect 5133 6747 5189 6803
rect 5964 6747 6020 6803
rect 6683 6747 6739 6803
rect 0 6205 8515 6666
rect 0 5565 8550 6142
rect 0 3987 8563 5469
rect 0 1414 8388 1866
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_0
timestamp 1763766357
transform 1 0 3194 0 1 3898
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_1
timestamp 1763766357
transform 1 0 2723 0 1 3898
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_2
timestamp 1763766357
transform 1 0 280 0 1 4038
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_3
timestamp 1763766357
transform 1 0 1064 0 1 4038
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_4
timestamp 1763766357
transform 1 0 4024 0 1 3755
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_5
timestamp 1763766357
transform 1 0 4181 0 1 3331
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_6
timestamp 1763766357
transform 1 0 750 0 1 3331
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_7
timestamp 1763766357
transform 1 0 593 0 1 3755
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_8
timestamp 1763766357
transform 1 0 3350 0 1 3614
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_9
timestamp 1763766357
transform 1 0 2566 0 1 3614
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_10
timestamp 1763766357
transform 1 0 3867 0 1 3473
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_11
timestamp 1763766357
transform 1 0 4337 0 1 3473
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_12
timestamp 1763766357
transform 1 0 2050 0 1 3473
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_13
timestamp 1763766357
transform 1 0 1579 0 1 3473
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_14
timestamp 1763766357
transform 1 0 1893 0 1 3331
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_15
timestamp 1763766357
transform 1 0 1736 0 1 3755
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_16
timestamp 1763766357
transform 1 0 4494 0 1 3614
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_17
timestamp 1763766357
transform 1 0 2207 0 1 4038
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_18
timestamp 1763766357
transform 1 0 1423 0 1 4038
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_19
timestamp 1763766357
transform 1 0 3710 0 1 3614
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_20
timestamp 1763766357
transform 1 0 907 0 1 3898
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_21
timestamp 1763766357
transform 1 0 436 0 1 3898
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_22
timestamp 1763766357
transform 1 0 2880 0 1 3755
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_23
timestamp 1763766357
transform 1 0 3037 0 1 3331
box -67 -48 67 47
use M1_POLY2_R270_256x8m81  M1_POLY2_R270_256x8m81_0
timestamp 1763766357
transform 0 -1 5126 -1 0 7063
box -48 -123 48 123
use M1_POLY24310591302019_256x8m81  M1_POLY24310591302019_256x8m81_0
timestamp 1763766357
transform 1 0 5600 0 1 7270
box -36 -80 36 78
use M1_POLY24310591302030_256x8m81  M1_POLY24310591302030_256x8m81_0
timestamp 1763766357
transform 1 0 6349 0 1 6653
box -95 -36 95 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_0
timestamp 1763766357
transform 1 0 5786 0 1 7043
box -36 -36 36 36
use M2_M1$$34864172_256x8m81  M2_M1$$34864172_256x8m81_0
timestamp 1763766357
transform -1 0 5103 0 1 7061
box -119 -46 119 46
use M2_M1$$34864172_256x8m81  M2_M1$$34864172_256x8m81_1
timestamp 1763766357
transform 0 1 5995 -1 0 6363
box -119 -46 119 46
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_0
timestamp 1763766357
transform 1 0 5623 0 1 7328
box -43 -122 43 122
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_1
timestamp 1763766357
transform 1 0 7160 0 1 6989
box -43 -122 43 122
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_2
timestamp 1763766357
transform 0 1 5989 -1 0 6874
box -43 -122 43 122
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_3
timestamp 1763766357
transform 0 1 6695 -1 0 6874
box -43 -122 43 122
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_4
timestamp 1763766357
transform 0 1 5077 -1 0 6880
box -43 -122 43 122
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_0
timestamp 1763766357
transform 1 0 6437 0 1 7363
box -44 -198 44 198
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_1
timestamp 1763766357
transform 1 0 5469 0 1 7403
box -44 -198 44 198
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_2
timestamp 1763766357
transform 1 0 5161 0 1 7403
box -44 -198 44 198
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_0
timestamp 1763766357
transform -1 0 8161 0 1 3335
box -44 -46 45 46
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_1
timestamp 1763766357
transform -1 0 7801 0 1 3759
box -44 -46 45 46
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_2
timestamp 1763766357
transform -1 0 5793 0 1 3618
box -44 -46 45 46
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_3
timestamp 1763766357
transform -1 0 6977 0 1 3477
box -44 -46 45 46
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_4
timestamp 1763766357
transform -1 0 6617 0 1 3900
box -44 -46 45 46
use M2_M1431059130200_256x8m81  M2_M1431059130200_256x8m81_0
timestamp 1763766357
transform 1 0 5747 0 1 7046
box -63 -34 63 34
use M3_M2$$43368492_256x8m81  M3_M2$$43368492_256x8m81_0
timestamp 1763766357
transform 0 1 5986 -1 0 6623
box -44 -123 44 123
use M3_M2$$43368492_256x8m81  M3_M2$$43368492_256x8m81_1
timestamp 1763766357
transform 0 1 6696 -1 0 6625
box -44 -123 44 123
use M3_M2$$43368492_256x8m81  M3_M2$$43368492_256x8m81_2
timestamp 1763766357
transform 0 1 5083 -1 0 7293
box -44 -123 44 123
use M3_M2$$43368492_256x8m81  M3_M2$$43368492_256x8m81_3
timestamp 1763766357
transform 0 1 5074 -1 0 6627
box -44 -123 44 123
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_0
timestamp 1763766357
transform 0 1 6590 -1 0 7210
box -45 -198 45 198
use nmos_1p2$$47342636_256x8m81  nmos_1p2$$47342636_256x8m81_0
timestamp 1763766357
transform 1 0 6341 0 1 7165
box -102 -44 130 170
use nmos_5p04310591302056_256x8m81  nmos_5p04310591302056_256x8m81_0
timestamp 1763766357
transform 1 0 5363 0 1 7168
box -88 -44 144 222
use nmos_5p04310591302056_256x8m81  nmos_5p04310591302056_256x8m81_1
timestamp 1763766357
transform 1 0 5203 0 1 7168
box -88 -44 144 222
use pmos_1p2$$47109164_256x8m81  pmos_1p2$$47109164_256x8m81_0
timestamp 1763766357
transform 1 0 6288 0 1 6733
box -216 -86 348 245
use xpredec1_bot_256x8m81  xpredec1_bot_256x8m81_0
timestamp 1763766357
transform 1 0 7155 0 1 562
box -74 852 1276 6007
use xpredec1_bot_256x8m81  xpredec1_bot_256x8m81_1
timestamp 1763766357
transform 1 0 4788 0 1 562
box -74 852 1276 6007
use xpredec1_bot_256x8m81  xpredec1_bot_256x8m81_2
timestamp 1763766357
transform 1 0 5971 0 1 562
box -74 852 1276 6007
use xpredec1_xa_256x8m81  xpredec1_xa_256x8m81_0
timestamp 1763766357
transform -1 0 3060 0 1 7450
box -46 -6036 774 228
use xpredec1_xa_256x8m81  xpredec1_xa_256x8m81_1
timestamp 1763766357
transform -1 0 4204 0 1 7450
box -46 -6036 774 228
use xpredec1_xa_256x8m81  xpredec1_xa_256x8m81_2
timestamp 1763766357
transform -1 0 1917 0 1 7450
box -46 -6036 774 228
use xpredec1_xa_256x8m81  xpredec1_xa_256x8m81_3
timestamp 1763766357
transform -1 0 773 0 1 7450
box -46 -6036 774 228
use xpredec1_xa_256x8m81  xpredec1_xa_256x8m81_4
timestamp 1763766357
transform 1 0 2874 0 1 7450
box -46 -6036 774 228
use xpredec1_xa_256x8m81  xpredec1_xa_256x8m81_5
timestamp 1763766357
transform 1 0 4018 0 1 7450
box -46 -6036 774 228
use xpredec1_xa_256x8m81  xpredec1_xa_256x8m81_6
timestamp 1763766357
transform 1 0 1731 0 1 7450
box -46 -6036 774 228
use xpredec1_xa_256x8m81  xpredec1_xa_256x8m81_7
timestamp 1763766357
transform 1 0 587 0 1 7450
box -46 -6036 774 228
<< labels >>
rlabel metal3 s 8399 4515 8399 4515 4 vdd
port 1 nsew
rlabel metal2 s 5029 7065 5029 7065 4 men
port 4 nsew
rlabel metal2 s 548 7632 548 7632 4 x[7]
port 5 nsew
rlabel metal2 s 796 7632 796 7632 4 x[6]
port 6 nsew
rlabel metal2 s 1692 7632 1692 7632 4 x[5]
port 7 nsew
rlabel metal2 s 1946 7632 1946 7632 4 x[4]
port 8 nsew
rlabel metal2 s 2834 7632 2834 7632 4 x[3]
port 9 nsew
rlabel metal2 s 3082 7632 3082 7632 4 x[2]
port 10 nsew
rlabel metal2 s 3997 7632 3997 7632 4 x[1]
port 11 nsew
rlabel metal2 s 4222 7632 4222 7632 4 x[0]
port 12 nsew
rlabel metal2 s 5623 7401 5623 7401 4 clk
port 15 nsew
rlabel metal2 s 5832 1695 5832 1695 4 A[2]
port 3 nsew
rlabel metal2 s 7016 1695 7016 1695 4 A[1]
port 13 nsew
rlabel metal2 s 8199 1695 8199 1695 4 A[0]
port 14 nsew
rlabel metal3 s 8269 1627 8269 1627 4 vss
port 2 nsew
rlabel metal3 s 8313 1488 8313 1488 4 vss
port 2 nsew
rlabel metal3 s 8399 5852 8399 5852 4 vss
port 2 nsew
rlabel metal3 s 8399 6449 8399 6449 4 vdd
port 1 nsew
rlabel metal3 s 8399 7179 8399 7179 4 vss
port 2 nsew
<< end >>
