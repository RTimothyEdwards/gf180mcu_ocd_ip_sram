magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< polysilicon >>
rect -1509 23 1509 36
rect -1509 -23 -1496 23
rect 1496 -23 1509 23
rect -1509 -36 1509 -23
<< polycontact >>
rect -1496 -23 1496 23
<< metal1 >>
rect -1504 23 1504 30
rect -1504 -23 -1496 23
rect 1496 -23 1504 23
rect -1504 -30 1504 -23
<< end >>
