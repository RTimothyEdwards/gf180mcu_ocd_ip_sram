magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< error_p >>
rect -75 0 -29 89
rect 85 0 131 89
<< nwell >>
rect -174 -86 230 175
<< pmos >>
rect 0 0 56 89
<< pdiff >>
rect -88 76 0 89
rect -88 13 -75 76
rect -29 13 0 76
rect -88 0 0 13
rect 56 76 144 89
rect 56 13 85 76
rect 131 13 144 76
rect 56 0 144 13
<< pdiffc >>
rect -75 13 -29 76
rect 85 13 131 76
<< polysilicon >>
rect 0 89 56 133
rect 0 -44 56 0
<< metal1 >>
rect -75 76 -29 89
rect -75 0 -29 13
rect 85 76 131 89
rect 85 0 131 13
<< labels >>
flabel pdiffc -40 44 -40 44 0 FreeSans 186 0 0 0 S
flabel pdiffc 96 44 96 44 0 FreeSans 186 0 0 0 D
<< end >>
