magic
tech gf180mcuD
magscale 1 10
timestamp 1763488735
<< nwell >>
rect 20780 64667 38804 64918
rect 20780 64635 27872 64667
rect 20780 64428 22995 64635
rect 24681 64429 27872 64635
rect 24682 64428 27872 64429
rect 31637 64617 38804 64667
rect 31637 64428 34834 64617
rect 36598 64428 38804 64617
<< psubdiff >>
rect 19420 23567 40130 23906
<< metal1 >>
rect 197 65044 60063 65744
rect 197 897 897 65044
rect 18028 64071 18537 65044
rect 19324 25153 20437 65044
rect 23958 64328 24509 65044
rect 28043 64328 28413 65044
rect 30616 64328 31194 65044
rect 35068 64198 35639 65044
rect 19170 24848 20437 25153
rect 38969 24848 40415 65044
rect 40953 64071 41462 65044
rect 19170 23900 19479 24848
rect 40106 23900 40415 24848
rect 59363 24557 60063 65044
rect 58864 24435 60063 24557
rect 19170 23573 40415 23900
rect 8934 1133 8989 1174
rect 9198 1133 9678 1188
rect 16457 1134 16822 1195
rect 18740 1022 19049 23122
rect 19170 1006 19479 23573
rect 34809 4069 35009 4101
rect 34974 3264 36262 3312
rect 40106 1006 40415 23573
rect 40536 1243 40845 23122
rect 58183 22092 58798 22144
rect 42864 1139 43376 1190
rect 42864 1138 43313 1139
rect 19170 897 40415 1006
rect 59363 897 60063 24435
rect 197 197 60063 897
<< metal2 >>
rect 197 65516 60063 65744
rect 494 64682 59766 65382
rect 494 197 1194 64682
rect 18029 18831 18537 64488
rect 18627 18986 18937 64682
rect 19170 64431 19479 64434
rect 19170 64292 20828 64431
rect 19170 63205 19479 64292
rect 20964 64198 21374 64682
rect 21538 64198 23021 64682
rect 24589 64198 25490 64682
rect 27267 64328 27732 64682
rect 34152 64198 34993 64682
rect 36558 64198 38047 64682
rect 38209 64198 38619 64682
rect 38759 64320 40161 64435
rect 19170 63066 20849 63205
rect 38759 63078 40161 63193
rect 19170 61993 19479 63066
rect 19170 61854 20849 61993
rect 38759 61866 40161 61981
rect 19170 60781 19479 61854
rect 19170 60642 20849 60781
rect 38759 60654 40161 60769
rect 19170 59569 19479 60642
rect 19170 59430 20849 59569
rect 38759 59442 40161 59557
rect 19170 58357 19479 59430
rect 19170 58218 20849 58357
rect 38759 58230 40161 58345
rect 19170 57145 19479 58218
rect 19170 57006 20849 57145
rect 38759 57018 40161 57133
rect 19170 55933 19479 57006
rect 19170 55794 20849 55933
rect 38759 55806 40161 55921
rect 19170 54721 19479 55794
rect 19170 54582 20849 54721
rect 38759 54594 40161 54709
rect 19170 53509 19479 54582
rect 19170 53370 20849 53509
rect 38759 53382 40161 53497
rect 19170 52297 19479 53370
rect 19170 52158 20849 52297
rect 38759 52170 40161 52285
rect 19170 51085 19479 52158
rect 19170 50946 20849 51085
rect 38759 50958 40161 51073
rect 19170 49873 19479 50946
rect 19170 49734 20849 49873
rect 38759 49746 40161 49861
rect 19170 48661 19479 49734
rect 19170 48522 20849 48661
rect 38759 48534 40161 48649
rect 19170 47449 19479 48522
rect 19170 47310 20849 47449
rect 38759 47322 40161 47437
rect 19170 46237 19479 47310
rect 19170 46098 20849 46237
rect 38759 46110 40161 46225
rect 19170 45025 19479 46098
rect 19170 44886 20849 45025
rect 38759 44898 40161 45013
rect 19170 43813 19479 44886
rect 19170 43674 20849 43813
rect 38759 43686 40161 43801
rect 19170 42601 19479 43674
rect 19170 42462 20849 42601
rect 38759 42474 40161 42589
rect 19170 41389 19479 42462
rect 19170 41250 20849 41389
rect 38759 41262 40161 41377
rect 19170 40177 19479 41250
rect 19170 40038 20849 40177
rect 38759 40050 40161 40165
rect 19170 38965 19479 40038
rect 19170 38826 20849 38965
rect 38759 38838 40161 38953
rect 19170 37753 19479 38826
rect 19170 37614 20849 37753
rect 38759 37626 40161 37741
rect 19170 36541 19479 37614
rect 19170 36402 20849 36541
rect 38759 36414 40161 36529
rect 19170 35329 19479 36402
rect 19170 35190 20849 35329
rect 38759 35202 40161 35317
rect 19170 34117 19479 35190
rect 19170 33978 20849 34117
rect 38759 33990 40161 34105
rect 19170 32905 19479 33978
rect 19170 32766 20849 32905
rect 38759 32778 40161 32893
rect 19170 31693 19479 32766
rect 19170 31554 20849 31693
rect 38759 31566 40161 31681
rect 19170 30481 19479 31554
rect 19170 30342 20849 30481
rect 38759 30354 40161 30469
rect 19170 29269 19479 30342
rect 19170 29130 20849 29269
rect 38759 29142 40161 29257
rect 19170 28057 19479 29130
rect 19170 27918 20849 28057
rect 38759 27930 40161 28045
rect 19170 26845 19479 27918
rect 19170 26706 20849 26845
rect 38759 26718 40161 26833
rect 19170 25633 19479 26706
rect 19170 25494 20849 25633
rect 38759 25506 40161 25621
rect 18803 18826 18897 18986
rect 17289 11644 17389 16713
rect 17480 11882 17580 16956
rect 17650 12121 17750 17198
rect 17826 12358 17926 17437
rect 18004 12596 18104 17973
rect 18178 12834 18278 18207
rect 18353 13072 18453 18460
rect 18544 13310 18644 18683
rect 1766 3293 1831 3524
rect 1304 3216 1831 3293
rect 2389 3402 2455 3517
rect 8443 3404 8509 3548
rect 2389 3359 2459 3402
rect 2389 3276 2517 3359
rect 2394 3275 2517 3276
rect 1304 3215 1797 3216
rect 1304 0 1461 3215
rect 1777 0 1934 1196
rect 2451 849 2517 3275
rect 8309 3338 8509 3404
rect 8309 945 8375 3338
rect 9055 3326 9120 3554
rect 8835 3261 9120 3326
rect 9537 3337 9602 3581
rect 10155 3428 10221 3579
rect 10155 3362 10316 3428
rect 9537 3280 9803 3337
rect 8835 1321 8900 3261
rect 8168 879 8375 945
rect 8643 1256 8900 1321
rect 8643 920 8708 1256
rect 2366 0 2522 849
rect 8168 840 8234 879
rect 8073 711 8234 840
rect 8636 834 8708 920
rect 8073 0 8229 711
rect 8544 0 8701 834
rect 8822 0 8979 1199
rect 9137 0 9294 1198
rect 9746 1085 9803 3280
rect 10250 1090 10316 3362
rect 16209 3287 16275 3545
rect 15595 3221 16275 3287
rect 16818 3293 16883 3523
rect 17139 3293 17200 3294
rect 9519 1028 9803 1085
rect 9519 832 9576 1028
rect 9992 1024 10316 1090
rect 9992 832 10058 1024
rect 9417 744 9576 832
rect 9417 0 9574 744
rect 9888 742 10058 832
rect 15596 826 15663 3221
rect 16818 3215 17200 3293
rect 9888 0 10045 742
rect 15595 0 15752 826
rect 16382 0 16539 1200
rect 16656 870 16813 876
rect 17139 870 17200 3215
rect 19170 2125 19479 25494
rect 25804 24709 26420 25314
rect 29030 24691 29185 24926
rect 27017 24531 29185 24691
rect 27017 24520 27171 24531
rect 22130 24359 27171 24520
rect 29295 24456 29450 24926
rect 22130 23003 22285 24359
rect 27353 24296 29450 24456
rect 27353 24278 27508 24296
rect 22379 24119 27508 24278
rect 29559 24222 29714 24926
rect 22379 23003 22534 24119
rect 27828 24061 29714 24222
rect 27828 23931 27983 24061
rect 29822 23986 29977 24918
rect 26810 23802 27983 23931
rect 26040 23771 27983 23802
rect 28074 23827 29977 23986
rect 26040 23643 26966 23771
rect 28074 23677 28229 23827
rect 30088 23752 30243 24926
rect 26040 23011 26196 23643
rect 27049 23568 28229 23677
rect 26289 23517 28229 23568
rect 28320 23592 30243 23752
rect 26289 23407 27204 23517
rect 28320 23442 28475 23592
rect 30351 23517 30506 24918
rect 31859 24748 32014 24926
rect 26289 23003 26444 23407
rect 27295 23282 28475 23442
rect 28566 23357 30506 23517
rect 31252 24588 32014 24748
rect 27295 23011 27450 23282
rect 28566 23196 28721 23357
rect 27544 23036 28721 23196
rect 31252 23162 31406 24588
rect 32123 24513 32278 24926
rect 31497 24353 32278 24513
rect 32387 24635 32543 24926
rect 32387 24476 32550 24635
rect 31497 23162 31653 24353
rect 32395 23162 32550 24476
rect 32652 24401 32807 24918
rect 32641 24240 32807 24401
rect 32641 23153 32796 24240
rect 32918 24044 33073 24918
rect 33181 24278 33336 24926
rect 33445 24513 33600 24926
rect 33709 24748 33865 24926
rect 33709 24588 35084 24748
rect 33445 24353 34838 24513
rect 33181 24119 33940 24278
rect 32918 23883 33694 24044
rect 33539 23153 33694 23883
rect 33785 23162 33940 24119
rect 34682 23162 34838 24353
rect 34928 23162 35084 24588
rect 34970 4074 35028 5910
rect 16656 809 17200 870
rect 16656 0 16813 809
rect 19555 0 19712 2026
rect 20304 1425 20394 2051
rect 20472 1761 20563 2051
rect 20472 1596 20950 1761
rect 20304 0 20461 1425
rect 20793 0 20950 1596
rect 21601 0 21758 4019
rect 22786 0 22943 4019
rect 23970 0 24126 4019
rect 28411 0 28568 1964
rect 35239 0 35396 4753
rect 36225 3298 36283 6575
rect 36157 3259 36283 3298
rect 37640 1931 38968 2088
rect 37640 0 37797 1931
rect 39046 1775 39137 2051
rect 38091 1619 39137 1775
rect 38091 0 38248 1619
rect 39216 1437 39306 2051
rect 38614 1280 39306 1437
rect 38614 0 38771 1280
rect 39385 0 39542 2269
rect 40106 2125 40415 23122
rect 40536 2125 40845 64682
rect 40953 18809 41461 64554
rect 59089 64018 59766 64682
rect 59088 23651 59766 64018
rect 42832 3293 42897 3526
rect 42451 3215 42897 3293
rect 43450 3359 43516 3515
rect 49509 3405 49566 3526
rect 43450 3275 43638 3359
rect 42451 871 42525 3215
rect 42451 797 42969 871
rect 42812 0 42969 797
rect 43280 0 43437 1191
rect 43572 941 43638 3275
rect 49435 3348 49566 3405
rect 43572 939 44012 941
rect 43572 875 44027 939
rect 43870 0 44027 875
rect 49435 849 49492 3348
rect 50117 3323 50175 3519
rect 49906 3267 50175 3323
rect 50648 3328 50713 3522
rect 50648 3271 50917 3328
rect 49906 849 49962 3267
rect 50299 2937 50305 2977
rect 50860 2937 50917 3271
rect 51266 3256 51332 3514
rect 57322 3279 57387 3555
rect 51266 3210 51468 3256
rect 51266 3190 51469 3210
rect 50859 1673 50916 2937
rect 50859 1612 50986 1673
rect 49376 0 49533 849
rect 49847 0 50004 849
rect 50126 0 50282 1202
rect 50641 0 50797 1200
rect 50929 849 50986 1612
rect 51405 849 51469 3190
rect 57174 3195 57387 3279
rect 57929 3281 57994 3521
rect 57929 3203 58397 3281
rect 57174 849 57240 3195
rect 50921 0 51077 849
rect 51392 0 51548 849
rect 57098 0 57255 849
rect 57686 0 57843 1199
rect 58240 1006 58397 3203
rect 58160 861 58397 1006
rect 58160 0 58317 861
rect 59066 197 59766 23651
<< metal3 >>
rect 1010 65516 1710 65942
rect 1868 65516 2568 65942
rect 2895 65516 3595 65942
rect 3753 65516 4453 65942
rect 4920 65516 5620 65942
rect 5778 65516 6478 65942
rect 6675 65516 7375 65942
rect 7533 65516 8233 65942
rect 8830 65516 9530 65942
rect 9688 65516 10388 65942
rect 10455 65516 11155 65942
rect 11313 65516 12013 65942
rect 12740 65516 13440 65942
rect 13598 65516 14298 65942
rect 14457 65516 15157 65942
rect 16090 65516 16790 65942
rect 16948 65516 17648 65942
rect 17760 65516 18460 65942
rect 18600 65516 19300 65942
rect 19663 65516 20363 65942
rect 20641 65516 21341 65942
rect 21497 65516 22197 65942
rect 22816 65516 23516 65942
rect 23966 65516 24666 65942
rect 24790 65516 25490 65942
rect 26013 65516 26713 65942
rect 27009 65516 27709 65942
rect 28067 65516 28767 65942
rect 28861 65516 29561 65942
rect 29851 65516 30551 65942
rect 30749 65516 31449 65942
rect 31548 65516 32248 65942
rect 32419 65516 33119 65942
rect 33276 65516 33976 65942
rect 34230 65516 34930 65942
rect 35475 65516 36175 65942
rect 36798 65516 37498 65942
rect 37983 65516 38683 65942
rect 39343 65516 40043 65942
rect 40282 65619 40982 65942
rect 41103 65619 41803 65942
rect 42103 65648 42803 65942
rect 42102 65516 42803 65648
rect 42961 65516 43661 65942
rect 44399 65516 45099 65942
rect 45256 65516 45956 65942
rect 46013 65516 46713 65942
rect 46871 65516 47571 65942
rect 48179 65516 48879 65942
rect 49036 65516 49736 65942
rect 49913 65516 50613 65942
rect 50771 65516 51471 65942
rect 51959 65516 52659 65942
rect 52816 65516 53516 65942
rect 53823 65516 54523 65942
rect 54681 65516 55381 65942
rect 55860 65516 56560 65942
rect 57163 65516 57863 65942
rect 58021 65516 58721 65942
rect 59066 65516 59766 65942
rect 42102 65515 42611 65516
rect 0 64682 60260 65382
rect 0 64116 709 64606
rect 19042 64291 19445 64432
rect 37782 64267 41389 64408
rect 0 63486 709 63976
rect 38000 63974 42103 64115
rect 59550 64093 60260 64582
rect 59550 63503 60260 63993
rect 0 62904 709 63394
rect 59550 62901 60260 63391
rect 0 62274 709 62764
rect 59550 62291 60260 62781
rect 0 61692 709 62182
rect 59550 61689 60260 62179
rect 0 61062 709 61552
rect 59550 61079 60260 61569
rect 0 60480 709 60970
rect 59550 60477 60260 60967
rect 0 59850 709 60340
rect 59550 59867 60260 60357
rect 0 59268 709 59758
rect 59550 59265 60260 59755
rect 0 58638 709 59128
rect 59550 58655 60260 59145
rect 0 58056 709 58546
rect 59550 58053 60260 58543
rect 0 57426 709 57916
rect 59550 57443 60260 57933
rect 0 56844 709 57334
rect 59550 56841 60260 57331
rect 0 56214 709 56704
rect 59550 56231 60260 56721
rect 0 55632 709 56122
rect 59550 55629 60260 56119
rect 0 55002 709 55492
rect 59550 55019 60260 55509
rect 0 54420 709 54910
rect 59550 54417 60260 54907
rect 0 53790 709 54280
rect 59550 53807 60260 54297
rect 0 53208 709 53698
rect 59550 53205 60260 53695
rect 0 52578 709 53068
rect 59550 52595 60260 53085
rect 0 51996 709 52486
rect 59550 51993 60260 52483
rect 0 51366 709 51856
rect 59550 51383 60260 51873
rect 0 50784 709 51274
rect 59550 50781 60260 51271
rect 0 50154 709 50644
rect 59550 50171 60260 50661
rect 0 49572 709 50062
rect 59550 49569 60260 50059
rect 0 48942 709 49432
rect 59550 48959 60260 49449
rect 0 48360 709 48850
rect 59550 48357 60260 48847
rect 0 47730 709 48220
rect 59550 47747 60260 48237
rect 0 47148 709 47638
rect 59550 47145 60260 47635
rect 0 46518 709 47008
rect 59550 46535 60260 47025
rect 0 45936 709 46426
rect 59550 45933 60260 46423
rect 0 45306 709 45796
rect 59550 45323 60260 45813
rect 0 44724 709 45214
rect 59550 44721 60260 45211
rect 0 44094 709 44584
rect 59550 44111 60260 44601
rect 0 43512 709 44002
rect 59550 43509 60260 43999
rect 0 42882 709 43372
rect 59550 42899 60260 43389
rect 0 42300 709 42790
rect 59550 42297 60260 42787
rect 0 41670 709 42160
rect 59550 41687 60260 42177
rect 0 41088 709 41578
rect 59550 41085 60260 41575
rect 0 40458 709 40948
rect 59550 40475 60260 40965
rect 0 39876 709 40366
rect 59550 39873 60260 40363
rect 0 39246 709 39736
rect 59550 39263 60260 39753
rect 0 38664 709 39154
rect 59550 38661 60260 39151
rect 0 38034 709 38524
rect 59550 38051 60260 38541
rect 0 37452 709 37942
rect 59550 37449 60260 37939
rect 0 36822 709 37312
rect 59550 36839 60260 37329
rect 0 36240 709 36730
rect 59550 36237 60260 36727
rect 0 35610 709 36100
rect 59550 35627 60260 36117
rect 0 35028 709 35493
rect 59550 35025 60260 35515
rect 0 34398 709 34888
rect 59550 34415 60260 34905
rect 0 33816 709 34306
rect 59550 33813 60260 34303
rect 0 33186 709 33676
rect 59550 33203 60260 33693
rect 0 32604 709 33094
rect 59550 32601 60260 33091
rect 0 31974 709 32464
rect 59550 31991 60260 32481
rect 0 31392 709 31882
rect 59550 31389 60260 31879
rect 0 30762 709 31252
rect 59550 30779 60260 31269
rect 0 30180 709 30670
rect 59550 30177 60260 30667
rect 0 29550 709 30040
rect 59550 29567 60260 30057
rect 0 28968 709 29458
rect 59550 28965 60260 29455
rect 0 28338 709 28828
rect 59550 28355 60260 28845
rect 0 27756 709 28246
rect 59550 27753 60260 28243
rect 0 27126 709 27616
rect 59550 27143 60260 27633
rect 0 26544 709 27034
rect 59551 27002 60260 27031
rect 59550 26541 60260 27002
rect 0 25914 709 26404
rect 59550 25931 60260 26421
rect 0 25332 709 25822
rect 59551 25780 60260 25819
rect 59550 25329 60260 25780
rect 0 24702 709 25192
rect 0 23834 709 24387
rect 17459 23968 19481 24170
rect 17529 23834 19481 23968
rect 0 20600 709 23546
rect 17529 22281 19049 23545
rect 25804 23407 26420 24803
rect 59550 24719 60260 25209
rect 40953 23834 42191 24170
rect 59550 23834 60260 24436
rect 19170 22276 20250 22943
rect 39294 22276 40415 22943
rect 40535 22279 42798 23545
rect 40535 22198 40845 22279
rect 18740 21699 20250 22198
rect 39294 21699 40845 22198
rect 17977 20969 20250 21605
rect 39328 20969 41466 21605
rect 16863 20615 20250 20798
rect 40534 20731 42942 20798
rect 16863 20600 20252 20615
rect 18740 20392 20252 20600
rect 39335 20600 42942 20731
rect 59550 20600 60260 23546
rect 0 18813 709 20200
rect 17186 19142 18249 20207
rect 18740 19297 20250 20392
rect 18740 19287 20247 19297
rect 39335 19196 40845 20600
rect 17186 18822 19479 19142
rect 40949 19129 43331 20194
rect 40106 18810 43331 19129
rect 59550 18813 60260 20200
rect 16965 18555 18683 18705
rect 16965 18319 18466 18470
rect 16965 18076 18289 18226
rect 16965 17835 18118 17986
rect 16963 17305 17940 17455
rect 16963 17060 17771 17210
rect 16963 16815 17606 16965
rect 19167 16827 20789 17304
rect 0 16115 709 16815
rect 16973 16569 17411 16720
rect 40540 16653 40854 16711
rect 18739 16630 40854 16653
rect 18739 16425 40853 16630
rect 16825 16115 43362 16425
rect 59550 16115 60260 16815
rect 18736 16114 43362 16115
rect 18736 16018 40853 16114
rect 18736 15934 19046 16018
rect 19170 15656 40376 15898
rect 0 14956 709 15656
rect 16825 15337 43362 15656
rect 19172 15262 39254 15337
rect 19172 15132 19482 15262
rect 40107 15225 40417 15337
rect 59551 15256 60260 15656
rect 59550 14956 60260 15256
rect 0 12620 709 14526
rect 16825 13637 42994 14176
rect 18538 13310 20582 13470
rect 39004 13310 41081 13470
rect 18345 13072 20582 13232
rect 39004 13072 41321 13232
rect 18174 12834 20582 12994
rect 39004 12834 41528 12994
rect 18001 12596 20582 12756
rect 39004 12596 41738 12756
rect 59550 12610 60260 14516
rect 0 10038 709 12420
rect 17821 12358 20582 12518
rect 39004 12358 41945 12518
rect 17642 12120 20582 12280
rect 39004 12120 42166 12280
rect 17483 11882 20582 12042
rect 39004 11882 42360 12042
rect 17282 11644 20582 11804
rect 39004 11644 42576 11804
rect 16877 10151 19479 11578
rect 39905 11407 42993 11510
rect 39905 11406 42994 11407
rect 38467 11354 42994 11406
rect 16877 10029 20636 10151
rect 38950 10136 42994 11354
rect 0 8434 709 9933
rect 16832 9052 19049 9924
rect 19170 9270 20636 10029
rect 40106 10033 42994 10136
rect 40106 9864 40428 10033
rect 59550 10028 60260 12410
rect 40246 9704 43638 9705
rect 40229 9421 43638 9704
rect 40229 9365 40914 9421
rect 16832 8712 20418 9052
rect 16832 8431 20636 8712
rect 18740 8289 20636 8431
rect 0 7132 709 8054
rect 16832 7122 19479 8044
rect 19679 7949 20636 8289
rect 38824 8671 40914 9365
rect 38824 8103 43638 8671
rect 59550 8424 60260 9923
rect 38824 7846 39780 8103
rect 40106 7702 43594 8042
rect 38902 7177 43594 7702
rect 40106 7122 43594 7177
rect 59550 7122 60260 8044
rect 16528 6958 20454 7020
rect 0 5715 709 6669
rect 16832 5706 20110 6660
rect 20393 6170 20454 6958
rect 38404 6958 43501 7020
rect 38404 6788 38466 6958
rect 36225 6726 38466 6788
rect 39058 6775 43220 6842
rect 36225 6519 36286 6726
rect 40536 6340 42899 6658
rect 20393 6108 29159 6170
rect 29097 5939 29159 6108
rect 29097 5877 35046 5939
rect 38832 5898 40415 6264
rect 18434 5455 20110 5706
rect 19724 5355 20110 5455
rect 0 4045 709 5326
rect 16537 4886 19479 5316
rect 19724 5114 20565 5355
rect 38836 5316 40415 5898
rect 40536 5386 43594 6340
rect 59550 5705 60260 6659
rect 19724 4961 20677 5114
rect 19724 4887 20679 4961
rect 38836 4888 43922 5316
rect 40455 4887 43922 4888
rect 16537 4413 20273 4811
rect 20356 4478 20679 4887
rect 39245 4413 43922 4810
rect 16580 4035 20622 4338
rect 38836 4035 43700 4338
rect 59550 4035 60260 5316
rect 0 2851 709 3949
rect 16580 3621 19049 3940
rect 40536 3621 43700 3940
rect 50835 3273 50913 3522
rect 40536 2855 43700 3173
rect 59550 2841 60260 3939
rect 40217 2651 42850 2652
rect 0 2006 709 2649
rect 40217 2405 43700 2651
rect 17006 2083 42931 2144
rect 59550 2006 60260 2299
rect 0 1760 60260 2006
rect 0 862 58933 1562
rect 59066 862 60260 1562
rect 494 0 1194 862
rect 1427 0 2127 862
rect 2409 0 3109 862
rect 3249 0 3949 311
rect 4089 0 4789 862
rect 4929 0 5629 862
rect 5769 0 6469 862
rect 6609 0 7309 311
rect 7449 0 8149 862
rect 8710 0 9410 862
rect 9969 0 10669 862
rect 10809 0 11509 311
rect 11649 0 12349 862
rect 12489 0 13189 862
rect 13329 0 14029 862
rect 14169 0 14869 311
rect 15337 0 16037 862
rect 16177 0 16877 862
rect 17087 0 17787 862
rect 17997 0 18697 862
rect 18907 0 19607 862
rect 19817 0 20517 862
rect 20727 0 21427 862
rect 21926 0 22626 311
rect 23115 0 23815 311
rect 24381 0 25081 311
rect 25221 0 25921 862
rect 26619 0 27319 311
rect 27459 0 28159 862
rect 28863 0 29563 311
rect 29703 0 30403 862
rect 30543 0 31243 311
rect 31383 0 32083 862
rect 32223 0 32923 311
rect 33063 0 33763 862
rect 33996 0 34696 862
rect 34913 0 35613 862
rect 35863 0 36563 311
rect 38120 0 38820 862
rect 39030 0 39730 862
rect 39940 0 40640 862
rect 40850 0 41550 862
rect 41760 0 42460 862
rect 42670 0 43370 862
rect 43606 0 44306 862
rect 44752 0 45452 311
rect 45592 0 46292 862
rect 46432 0 47132 862
rect 47272 0 47972 862
rect 48112 0 48812 311
rect 48952 0 49652 862
rect 50211 0 50911 862
rect 51472 0 52172 862
rect 52312 0 53012 311
rect 53152 0 53852 862
rect 53992 0 54692 862
rect 54832 0 55532 862
rect 55672 0 56372 311
rect 56712 0 57412 862
rect 57693 0 58393 862
rect 59066 0 59766 862
use 512x8M8W_PWR_512x8m81  512x8M8W_PWR_512x8m81_0
timestamp 1763482574
transform 1 0 0 0 1 -341
box 1338 4614 58383 24803
use control_512x8_512x8m81  control_512x8_512x8m81_0
timestamp 1763486358
transform 1 0 19273 0 1 2956
box -2537 -1052 22252 21087
use G_ring_512x8m81  G_ring_512x8m81_0
timestamp 1763482574
transform 1 0 197 0 1 -341
box 0 341 59871 65718
use GF018_512x8M8WM1_lef_512x8m81  GF018_512x8M8WM1_lef_512x8m81_0
timestamp 1763482574
transform 1 0 0 0 1 -341
box 0 341 60260 66283
use lcol4_512_512x8m81  lcol4_512_512x8m81_0
timestamp 1763486358
transform 1 0 2044 0 1 3172
box -830 -2043 15967 61786
use M1_PSUB4310591302010_512x8m81  M1_PSUB4310591302010_512x8m81_0
timestamp 1763476864
transform 1 0 37597 0 1 1605
box -2018 -800 2018 800
use M1_PSUB4310591302014_512x8m81  M1_PSUB4310591302014_512x8m81_0
timestamp 1763476864
transform 1 0 24082 0 1 1605
box -4048 -800 4048 800
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_0
timestamp 1763476864
transform 1 0 39671 0 1 25564
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_1
timestamp 1763476864
transform 1 0 39671 0 1 26776
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_2
timestamp 1763476864
transform 1 0 39671 0 1 27989
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_3
timestamp 1763476864
transform 1 0 39671 0 1 29200
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_4
timestamp 1763476864
transform 1 0 39671 0 1 30412
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_5
timestamp 1763476864
transform 1 0 39671 0 1 31624
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_6
timestamp 1763476864
transform 1 0 39671 0 1 32836
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_7
timestamp 1763476864
transform 1 0 19914 0 1 32837
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_8
timestamp 1763476864
transform 1 0 19914 0 1 31624
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_9
timestamp 1763476864
transform 1 0 19914 0 1 30412
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_10
timestamp 1763476864
transform 1 0 19914 0 1 29200
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_11
timestamp 1763476864
transform 1 0 19914 0 1 25567
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_12
timestamp 1763476864
transform 1 0 19914 0 1 26777
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_13
timestamp 1763476864
transform 1 0 19914 0 1 27987
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_14
timestamp 1763476864
transform 1 0 19914 0 1 63136
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_15
timestamp 1763476864
transform 1 0 19914 0 1 61924
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_16
timestamp 1763476864
transform 1 0 19914 0 1 60712
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_17
timestamp 1763476864
transform 1 0 19914 0 1 59500
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_18
timestamp 1763476864
transform 1 0 19914 0 1 58288
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_19
timestamp 1763476864
transform 1 0 19914 0 1 57076
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_20
timestamp 1763476864
transform 1 0 19914 0 1 55864
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_21
timestamp 1763476864
transform 1 0 19914 0 1 54652
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_22
timestamp 1763476864
transform 1 0 19914 0 1 53440
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_23
timestamp 1763476864
transform 1 0 19914 0 1 52228
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_24
timestamp 1763476864
transform 1 0 19914 0 1 51016
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_25
timestamp 1763476864
transform 1 0 19914 0 1 49804
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_26
timestamp 1763476864
transform 1 0 19914 0 1 48592
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_27
timestamp 1763476864
transform 1 0 19914 0 1 47380
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_28
timestamp 1763476864
transform 1 0 19914 0 1 46168
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_29
timestamp 1763476864
transform 1 0 19914 0 1 44956
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_30
timestamp 1763476864
transform 1 0 19914 0 1 43744
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_31
timestamp 1763476864
transform 1 0 19914 0 1 42532
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_32
timestamp 1763476864
transform 1 0 19914 0 1 41320
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_33
timestamp 1763476864
transform 1 0 19914 0 1 40108
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_34
timestamp 1763476864
transform 1 0 19914 0 1 38896
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_35
timestamp 1763476864
transform 1 0 19914 0 1 37684
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_36
timestamp 1763476864
transform 1 0 19914 0 1 36472
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_37
timestamp 1763476864
transform 1 0 19914 0 1 35260
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_38
timestamp 1763476864
transform 1 0 19914 0 1 34048
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_39
timestamp 1763476864
transform 1 0 19914 0 1 64348
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_40
timestamp 1763476864
transform 1 0 39671 0 1 59500
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_41
timestamp 1763476864
transform 1 0 39671 0 1 60712
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_42
timestamp 1763476864
transform 1 0 39671 0 1 61925
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_43
timestamp 1763476864
transform 1 0 39671 0 1 63136
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_44
timestamp 1763476864
transform 1 0 39671 0 1 64376
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_45
timestamp 1763476864
transform 1 0 39671 0 1 34048
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_46
timestamp 1763476864
transform 1 0 39671 0 1 35260
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_47
timestamp 1763476864
transform 1 0 39671 0 1 36472
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_48
timestamp 1763476864
transform 1 0 39671 0 1 37684
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_49
timestamp 1763476864
transform 1 0 39671 0 1 38896
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_50
timestamp 1763476864
transform 1 0 39671 0 1 40108
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_51
timestamp 1763476864
transform 1 0 39671 0 1 41320
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_52
timestamp 1763476864
transform 1 0 39671 0 1 42532
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_53
timestamp 1763476864
transform 1 0 39671 0 1 43744
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_54
timestamp 1763476864
transform 1 0 39671 0 1 44956
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_55
timestamp 1763476864
transform 1 0 39671 0 1 46168
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_56
timestamp 1763476864
transform 1 0 39671 0 1 47380
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_57
timestamp 1763476864
transform 1 0 39671 0 1 48592
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_58
timestamp 1763476864
transform 1 0 39671 0 1 49804
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_59
timestamp 1763476864
transform 1 0 39671 0 1 51016
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_60
timestamp 1763476864
transform 1 0 39671 0 1 52228
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_61
timestamp 1763476864
transform 1 0 39671 0 1 53439
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_62
timestamp 1763476864
transform 1 0 39671 0 1 54672
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_63
timestamp 1763476864
transform 1 0 39671 0 1 55864
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_64
timestamp 1763476864
transform 1 0 39671 0 1 57076
box -487 -46 487 46
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_65
timestamp 1763476864
transform 1 0 39671 0 1 58288
box -487 -46 487 46
use M2_M1$$201260076_512x8m81  M2_M1$$201260076_512x8m81_0
timestamp 1763476864
transform -1 0 40260 0 1 13217
box -119 -9872 119 9872
use M2_M1$$201260076_512x8m81  M2_M1$$201260076_512x8m81_1
timestamp 1763476864
transform -1 0 40691 0 1 13217
box -119 -9872 119 9872
use M2_M1$$201260076_512x8m81  M2_M1$$201260076_512x8m81_2
timestamp 1763476864
transform 1 0 19325 0 1 13217
box -119 -9872 119 9872
use M2_M1$$201260076_512x8m81  M2_M1$$201260076_512x8m81_3
timestamp 1763476864
transform 1 0 18895 0 1 13217
box -119 -9872 119 9872
use M2_M1$$201261100_512x8m81  M2_M1$$201261100_512x8m81_0
timestamp 1763476864
transform -1 0 40691 0 1 2547
box -119 -351 119 351
use M2_M1$$201261100_512x8m81  M2_M1$$201261100_512x8m81_1
timestamp 1763476864
transform -1 0 40260 0 1 2547
box -119 -351 119 351
use M2_M1$$201261100_512x8m81  M2_M1$$201261100_512x8m81_2
timestamp 1763476864
transform 1 0 19325 0 1 2547
box -119 -351 119 351
use M2_M1$$201261100_512x8m81  M2_M1$$201261100_512x8m81_3
timestamp 1763476864
transform 1 0 18895 0 1 2547
box -119 -351 119 351
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_0
timestamp 1763476864
transform 1 0 43359 0 1 1154
box -63 -34 63 34
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_1
timestamp 1763476864
transform 1 0 34990 0 1 4085
box -63 -34 63 34
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_2
timestamp 1763476864
transform 1 0 57765 0 1 1164
box -63 -34 63 34
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_3
timestamp 1763476864
transform 1 0 36212 0 1 3280
box -63 -34 63 34
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_4
timestamp 1763476864
transform 1 0 50720 0 1 1163
box -63 -34 63 34
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_5
timestamp 1763476864
transform 1 0 50205 0 1 1163
box -63 -34 63 34
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_6
timestamp 1763476864
transform 1 0 16461 0 1 1164
box -63 -34 63 34
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_7
timestamp 1763476864
transform 1 0 9246 0 1 1164
box -63 -34 63 34
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_8
timestamp 1763476864
transform 1 0 8901 0 1 1164
box -63 -34 63 34
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_9
timestamp 1763476864
transform 1 0 1856 0 1 1163
box -63 -34 63 34
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_10
timestamp 1763476864
transform 1 0 28490 0 1 1938
box -63 -34 63 34
use M2_M1431059130203_512x8m81  M2_M1431059130203_512x8m81_0
timestamp 1763476864
transform 1 0 18271 0 1 24002
box -200 -156 200 156
use M2_M1431059130204_512x8m81  M2_M1431059130204_512x8m81_0
timestamp 1763476864
transform 1 0 18293 0 1 64365
box -200 -113 200 113
use M2_M1431059130204_512x8m81  M2_M1431059130204_512x8m81_1
timestamp 1763476864
transform 1 0 41198 0 1 64435
box -200 -113 200 113
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_0
timestamp 1763476864
transform 1 0 41870 0 1 24456
box -34 -63 34 63
use M2_M14310591302012_512x8m81  M2_M14310591302012_512x8m81_0
timestamp 1763476864
transform 1 0 19319 0 1 24003
box -113 -156 113 156
use m2m3_512x8m81  m2m3_512x8m81_0
timestamp 1763482574
transform 1 0 41027 0 1 11644
box -75 0 2478 7071
use M3_M2$$201248812_512x8m81  M3_M2$$201248812_512x8m81_0
timestamp 1763476864
transform -1 0 40691 0 1 8917
box -119 -732 119 732
use M3_M2$$201248812_512x8m81  M3_M2$$201248812_512x8m81_1
timestamp 1763476864
transform -1 0 40260 0 1 10628
box -119 -732 119 732
use M3_M2$$201248812_512x8m81  M3_M2$$201248812_512x8m81_2
timestamp 1763476864
transform 1 0 19325 0 1 10823
box -119 -732 119 732
use M3_M2$$201248812_512x8m81  M3_M2$$201248812_512x8m81_3
timestamp 1763476864
transform 1 0 18895 0 1 9177
box -119 -732 119 732
use M3_M2$$201249836_512x8m81  M3_M2$$201249836_512x8m81_0
timestamp 1763483012
transform -1 0 40260 0 1 7582
box -119 -427 119 427
use M3_M2$$201249836_512x8m81  M3_M2$$201249836_512x8m81_1
timestamp 1763483012
transform -1 0 40691 0 1 5863
box -119 -427 119 427
use M3_M2$$201249836_512x8m81  M3_M2$$201249836_512x8m81_2
timestamp 1763483012
transform 1 0 19325 0 1 7582
box -119 -427 119 427
use M3_M2$$201249836_512x8m81  M3_M2$$201249836_512x8m81_3
timestamp 1763483012
transform 1 0 18895 0 1 5913
box -119 -427 119 427
use M3_M2$$201250860_512x8m81  M3_M2$$201250860_512x8m81_0
timestamp 1763476864
transform -1 0 39553 0 1 4612
box -266 -198 266 198
use M3_M2$$201250860_512x8m81  M3_M2$$201250860_512x8m81_1
timestamp 1763476864
transform 1 0 20002 0 1 4612
box -266 -198 266 198
use M3_M2$$201251884_512x8m81  M3_M2$$201251884_512x8m81_0
timestamp 1763476864
transform 1 0 26112 0 1 24756
box -266 -46 266 46
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_0
timestamp 1763476864
transform 1 0 20180 0 1 2522
box -45 -122 45 123
use M3_M2$$201253932_512x8m81  M3_M2$$201253932_512x8m81_0
timestamp 1763476864
transform 1 0 40260 0 1 5712
box -119 -808 119 511
use M3_M2$$201254956_512x8m81  M3_M2$$201254956_512x8m81_0
timestamp 1763476864
transform 1 0 19325 0 1 9636
box -119 -351 119 351
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_0
timestamp 1763476864
transform 1 0 19914 0 1 34048
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_1
timestamp 1763476864
transform 1 0 39671 0 1 26776
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_2
timestamp 1763476864
transform 1 0 39671 0 1 27989
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_3
timestamp 1763476864
transform 1 0 39671 0 1 29200
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_4
timestamp 1763476864
transform 1 0 39671 0 1 30412
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_5
timestamp 1763476864
transform 1 0 39671 0 1 31624
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_6
timestamp 1763476864
transform 1 0 39671 0 1 32836
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_7
timestamp 1763476864
transform 1 0 19914 0 1 32836
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_8
timestamp 1763476864
transform 1 0 19914 0 1 31624
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_9
timestamp 1763476864
transform 1 0 19914 0 1 30412
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_10
timestamp 1763476864
transform 1 0 19914 0 1 29200
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_11
timestamp 1763476864
transform 1 0 19914 0 1 27987
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_12
timestamp 1763476864
transform 1 0 19914 0 1 26779
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_13
timestamp 1763476864
transform 1 0 19914 0 1 25567
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_14
timestamp 1763476864
transform 1 0 19914 0 1 55864
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_15
timestamp 1763476864
transform 1 0 19914 0 1 54652
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_16
timestamp 1763476864
transform 1 0 19914 0 1 53440
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_17
timestamp 1763476864
transform 1 0 19914 0 1 52228
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_18
timestamp 1763476864
transform 1 0 19914 0 1 51016
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_19
timestamp 1763476864
transform 1 0 19914 0 1 49804
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_20
timestamp 1763476864
transform 1 0 19914 0 1 48592
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_21
timestamp 1763476864
transform 1 0 19914 0 1 47380
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_22
timestamp 1763476864
transform 1 0 19914 0 1 46168
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_23
timestamp 1763476864
transform 1 0 19914 0 1 44956
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_24
timestamp 1763476864
transform 1 0 19914 0 1 43744
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_25
timestamp 1763476864
transform 1 0 19914 0 1 42532
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_26
timestamp 1763476864
transform 1 0 19914 0 1 41320
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_27
timestamp 1763476864
transform 1 0 19914 0 1 40108
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_28
timestamp 1763476864
transform 1 0 19914 0 1 38896
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_29
timestamp 1763476864
transform 1 0 19914 0 1 37684
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_30
timestamp 1763476864
transform 1 0 19914 0 1 36472
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_31
timestamp 1763476864
transform 1 0 19914 0 1 35260
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_32
timestamp 1763476864
transform 1 0 19914 0 1 34048
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_33
timestamp 1763476864
transform 1 0 19914 0 1 64348
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_34
timestamp 1763476864
transform 1 0 19914 0 1 63136
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_35
timestamp 1763476864
transform 1 0 19914 0 1 61924
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_36
timestamp 1763476864
transform 1 0 19914 0 1 60712
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_37
timestamp 1763476864
transform 1 0 19914 0 1 59500
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_38
timestamp 1763476864
transform 1 0 19914 0 1 58288
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_39
timestamp 1763476864
transform 1 0 19914 0 1 57076
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_40
timestamp 1763476864
transform 1 0 39671 0 1 34048
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_41
timestamp 1763476864
transform 1 0 39671 0 1 35260
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_42
timestamp 1763476864
transform 1 0 39671 0 1 36472
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_43
timestamp 1763476864
transform 1 0 39671 0 1 37684
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_44
timestamp 1763476864
transform 1 0 39671 0 1 38896
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_45
timestamp 1763476864
transform 1 0 39671 0 1 40108
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_46
timestamp 1763476864
transform 1 0 39671 0 1 41320
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_47
timestamp 1763476864
transform 1 0 39671 0 1 42532
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_48
timestamp 1763476864
transform 1 0 39671 0 1 43744
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_49
timestamp 1763476864
transform 1 0 39671 0 1 44956
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_50
timestamp 1763476864
transform 1 0 39671 0 1 46168
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_51
timestamp 1763476864
transform 1 0 39671 0 1 47380
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_52
timestamp 1763476864
transform 1 0 39671 0 1 48592
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_53
timestamp 1763476864
transform 1 0 39671 0 1 49804
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_54
timestamp 1763476864
transform 1 0 39671 0 1 51016
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_55
timestamp 1763476864
transform 1 0 39671 0 1 52228
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_56
timestamp 1763476864
transform 1 0 39671 0 1 53439
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_57
timestamp 1763476864
transform 1 0 39671 0 1 54672
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_58
timestamp 1763476864
transform 1 0 39671 0 1 55864
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_59
timestamp 1763476864
transform 1 0 39671 0 1 57076
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_60
timestamp 1763476864
transform 1 0 39671 0 1 58288
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_61
timestamp 1763476864
transform 1 0 39671 0 1 59500
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_62
timestamp 1763476864
transform 1 0 39671 0 1 60712
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_63
timestamp 1763476864
transform 1 0 39671 0 1 61925
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_64
timestamp 1763476864
transform 1 0 39671 0 1 63136
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_65
timestamp 1763476864
transform 1 0 39671 0 1 64376
box -487 -46 487 46
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_66
timestamp 1763476864
transform 1 0 39671 0 1 25564
box -487 -46 487 46
use M3_M2$$201412652_512x8m81  M3_M2$$201412652_512x8m81_0
timestamp 1763476864
transform -1 0 40260 0 1 21286
box -119 -275 119 275
use M3_M2$$201412652_512x8m81  M3_M2$$201412652_512x8m81_1
timestamp 1763476864
transform -1 0 40260 0 1 22609
box -119 -275 119 275
use M3_M2$$201412652_512x8m81  M3_M2$$201412652_512x8m81_2
timestamp 1763476864
transform 1 0 19325 0 1 22609
box -119 -275 119 275
use M3_M2$$201412652_512x8m81  M3_M2$$201412652_512x8m81_3
timestamp 1763476864
transform 1 0 19325 0 1 21286
box -119 -275 119 275
use M3_M2$$201413676_512x8m81  M3_M2$$201413676_512x8m81_0
timestamp 1763476864
transform -1 0 40691 0 1 21948
box -119 -198 119 198
use M3_M2$$201413676_512x8m81  M3_M2$$201413676_512x8m81_1
timestamp 1763476864
transform 1 0 18895 0 1 21948
box -119 -198 119 198
use M3_M2$$201413676_512x8m81  M3_M2$$201413676_512x8m81_2
timestamp 1763476864
transform 1 0 19325 0 1 5101
box -119 -198 119 198
use M3_M2$$201414700_512x8m81  M3_M2$$201414700_512x8m81_0
timestamp 1763476864
transform -1 0 40691 0 1 22913
box -119 -579 119 579
use M3_M2$$201414700_512x8m81  M3_M2$$201414700_512x8m81_1
timestamp 1763476864
transform 1 0 18895 0 1 22913
box -119 -579 119 579
use M3_M2$$201415724_512x8m81  M3_M2$$201415724_512x8m81_0
timestamp 1763476864
transform -1 0 40691 0 1 19779
box -119 -584 119 884
use M3_M2$$201415724_512x8m81  M3_M2$$201415724_512x8m81_1
timestamp 1763476864
transform 1 0 18895 0 1 19879
box -119 -584 119 884
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_0
timestamp 1763476864
transform -1 0 40260 0 1 2529
box -119 -123 119 123
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_1
timestamp 1763476864
transform -1 0 40691 0 1 3780
box -119 -123 119 123
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_2
timestamp 1763476864
transform -1 0 40260 0 1 4187
box -119 -123 119 123
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_3
timestamp 1763476864
transform -1 0 40691 0 1 3032
box -119 -123 119 123
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_4
timestamp 1763476864
transform -1 0 40260 0 1 18969
box -119 -123 119 123
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_5
timestamp 1763476864
transform 1 0 19325 0 1 2520
box -119 -123 119 123
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_6
timestamp 1763476864
transform 1 0 18895 0 1 3003
box -119 -123 119 123
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_7
timestamp 1763476864
transform 1 0 19325 0 1 4187
box -119 -123 119 123
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_8
timestamp 1763476864
transform 1 0 18895 0 1 3780
box -119 -123 119 123
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_9
timestamp 1763476864
transform 1 0 19325 0 1 18982
box -119 -123 119 123
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_10
timestamp 1763476864
transform 1 0 19325 0 1 17082
box -119 -123 119 123
use M3_M2431059130201_512x8m81  M3_M2431059130201_512x8m81_0
timestamp 1763476864
transform 0 -1 34983 1 0 5906
box -35 -63 35 63
use M3_M2431059130201_512x8m81  M3_M2431059130201_512x8m81_1
timestamp 1763476864
transform 1 0 36255 0 1 6582
box -35 -63 35 63
use M3_M2431059130202_512x8m81  M3_M2431059130202_512x8m81_0
timestamp 1763476864
transform 1 0 18271 0 1 24003
box -200 -156 200 156
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_0
timestamp 1763476864
transform 1 0 40689 0 1 14002
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_1
timestamp 1763476864
transform 1 0 40689 0 1 13761
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_2
timestamp 1763476864
transform 1 0 17352 0 1 11724
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_3
timestamp 1763476864
transform 1 0 17527 0 1 16889
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_4
timestamp 1763476864
transform 1 0 17546 0 1 11962
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_5
timestamp 1763476864
transform 1 0 17696 0 1 17134
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_6
timestamp 1763476864
transform 1 0 17715 0 1 12186
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_7
timestamp 1763476864
transform 1 0 17872 0 1 17378
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_8
timestamp 1763476864
transform 1 0 17891 0 1 12448
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_9
timestamp 1763476864
transform 1 0 18050 0 1 17912
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_10
timestamp 1763476864
transform 1 0 18069 0 1 12681
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_11
timestamp 1763476864
transform 1 0 18225 0 1 18146
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_12
timestamp 1763476864
transform 1 0 18245 0 1 12921
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_13
timestamp 1763476864
transform 1 0 18400 0 1 18389
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_14
timestamp 1763476864
transform 1 0 18420 0 1 13145
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_15
timestamp 1763476864
transform 1 0 18611 0 1 18623
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_16
timestamp 1763476864
transform 1 0 18611 0 1 13387
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_17
timestamp 1763476864
transform 1 0 18902 0 1 14002
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_18
timestamp 1763476864
transform 1 0 18902 0 1 13761
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_19
timestamp 1763476864
transform 1 0 17335 0 1 16644
box -63 -63 63 63
use M3_M2431059130206_512x8m81  M3_M2431059130206_512x8m81_0
timestamp 1763476864
transform 1 0 19319 0 1 24003
box -113 -156 113 156
use M3_M2431059130207_512x8m81  M3_M2431059130207_512x8m81_0
timestamp 1763476864
transform 1 0 30716 0 1 2114
box -63 -35 63 35
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_0
timestamp 1763476864
transform 1 0 41204 0 1 21461
box -200 -113 200 113
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_1
timestamp 1763476864
transform 1 0 41204 0 1 21149
box -200 -113 200 113
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_2
timestamp 1763476864
transform 1 0 18271 0 1 21426
box -200 -113 200 113
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_3
timestamp 1763476864
transform 1 0 18271 0 1 21107
box -200 -113 200 113
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_4
timestamp 1763476864
transform 1 0 18293 0 1 64365
box -200 -113 200 113
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_5
timestamp 1763476864
transform 1 0 41198 0 1 64435
box -200 -113 200 113
use M3_M24310591302011_512x8m81  M3_M24310591302011_512x8m81_0
timestamp 1763476864
transform 1 0 41207 0 1 24003
box -243 -156 243 156
use M3_M24310591302013_512x8m81  M3_M24310591302013_512x8m81_0
timestamp 1763476864
transform 1 0 40688 0 1 16360
box -99 -317 99 317
use M3_M24310591302013_512x8m81  M3_M24310591302013_512x8m81_1
timestamp 1763476864
transform 1 0 40246 0 1 15564
box -99 -317 99 317
use M3_M24310591302013_512x8m81  M3_M24310591302013_512x8m81_2
timestamp 1763476864
transform 1 0 18893 0 1 16300
box -99 -317 99 317
use M3_M24310591302013_512x8m81  M3_M24310591302013_512x8m81_3
timestamp 1763476864
transform 1 0 19324 0 1 15503
box -99 -317 99 317
use M3_M24310591302015_512x8m81  M3_M24310591302015_512x8m81_0
timestamp 1763476864
transform 1 0 41194 0 1 19538
box -200 -634 200 634
use M3_M24310591302015_512x8m81  M3_M24310591302015_512x8m81_1
timestamp 1763476864
transform 1 0 18276 0 1 19513
box -200 -634 200 634
use power_a_512x8m81  power_a_512x8m81_0
timestamp 1763476864
transform -1 0 48812 0 1 197
box 0 -197 700 700
use power_a_512x8m81  power_a_512x8m81_1
timestamp 1763476864
transform -1 0 56372 0 1 197
box 0 -197 700 700
use power_a_512x8m81  power_a_512x8m81_2
timestamp 1763476864
transform 1 0 52312 0 1 197
box 0 -197 700 700
use power_a_512x8m81  power_a_512x8m81_3
timestamp 1763476864
transform 1 0 32223 0 1 197
box 0 -197 700 700
use power_a_512x8m81  power_a_512x8m81_4
timestamp 1763476864
transform 1 0 36734 0 1 197
box 0 -197 700 700
use power_a_512x8m81  power_a_512x8m81_5
timestamp 1763476864
transform 1 0 30543 0 1 197
box 0 -197 700 700
use power_a_512x8m81  power_a_512x8m81_6
timestamp 1763476864
transform 1 0 35863 0 1 197
box 0 -197 700 700
use power_a_512x8m81  power_a_512x8m81_7
timestamp 1763476864
transform 1 0 44752 0 1 197
box 0 -197 700 700
use power_a_512x8m81  power_a_512x8m81_8
timestamp 1763476864
transform -1 0 23815 0 1 197
box 0 -197 700 700
use power_a_512x8m81  power_a_512x8m81_9
timestamp 1763476864
transform -1 0 22626 0 1 197
box 0 -197 700 700
use power_a_512x8m81  power_a_512x8m81_10
timestamp 1763476864
transform -1 0 7309 0 1 197
box 0 -197 700 700
use power_a_512x8m81  power_a_512x8m81_11
timestamp 1763476864
transform -1 0 14869 0 1 197
box 0 -197 700 700
use power_a_512x8m81  power_a_512x8m81_12
timestamp 1763476864
transform 1 0 28863 0 1 197
box 0 -197 700 700
use power_a_512x8m81  power_a_512x8m81_13
timestamp 1763476864
transform 1 0 10809 0 1 197
box 0 -197 700 700
use power_a_512x8m81  power_a_512x8m81_14
timestamp 1763476864
transform 1 0 24381 0 1 197
box 0 -197 700 700
use power_a_512x8m81  power_a_512x8m81_15
timestamp 1763476864
transform 1 0 3249 0 1 197
box 0 -197 700 700
use power_a_512x8m81  power_a_512x8m81_16
timestamp 1763476864
transform 1 0 26619 0 1 197
box 0 -197 700 700
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_0
timestamp 1763476864
transform 1 0 10813 0 1 64241
box -357 441 1199 1701
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_1
timestamp 1763476864
transform 1 0 7033 0 1 64241
box -357 441 1199 1701
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_2
timestamp 1763476864
transform 1 0 3253 0 1 64241
box -357 441 1199 1701
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_3
timestamp 1763476864
transform 1 0 52316 0 1 64241
box -357 441 1199 1701
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_4
timestamp 1763476864
transform 1 0 48536 0 1 64241
box -357 441 1199 1701
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_5
timestamp 1763476864
transform 1 0 44756 0 1 64241
box -357 441 1199 1701
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_6
timestamp 1763476864
transform 1 0 32776 0 1 64241
box -357 441 1199 1701
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_0
timestamp 1763476864
transform -1 0 29203 0 1 64241
box -357 441 342 1701
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_1
timestamp 1763476864
transform -1 0 27351 0 1 64241
box -357 441 342 1701
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_2
timestamp 1763476864
transform -1 0 25132 0 1 64241
box -357 441 342 1701
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_3
timestamp 1763476864
transform -1 0 21839 0 1 64241
box -357 441 342 1701
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_4
timestamp 1763476864
transform -1 0 18942 0 1 64241
box -357 441 342 1701
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_5
timestamp 1763476864
transform -1 0 14799 0 1 64241
box -357 441 342 1701
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_6
timestamp 1763476864
transform -1 0 56202 0 1 64241
box -357 441 342 1701
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_7
timestamp 1763476864
transform -1 0 40625 0 1 64241
box -357 441 342 1701
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_8
timestamp 1763476864
transform -1 0 59408 0 1 64241
box -357 441 342 1701
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_9
timestamp 1763476864
transform -1 0 38325 0 1 64241
box -357 441 342 1701
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_10
timestamp 1763476864
transform -1 0 34573 0 1 64241
box -357 441 342 1701
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_11
timestamp 1763476864
transform -1 0 31890 0 1 64241
box -357 441 342 1701
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_12
timestamp 1763476864
transform -1 0 37140 0 1 64241
box -357 441 342 1701
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_0
timestamp 1763476864
transform -1 0 18810 0 1 64241
box 349 1275 1049 1701
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_1
timestamp 1763476864
transform -1 0 29117 0 1 64241
box 349 1275 1049 1701
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_2
timestamp 1763476864
transform -1 0 27063 0 1 64241
box 349 1275 1049 1701
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_3
timestamp 1763476864
transform -1 0 25016 0 1 64241
box 349 1275 1049 1701
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_4
timestamp 1763476864
transform -1 0 23866 0 1 64241
box 349 1275 1049 1701
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_5
timestamp 1763476864
transform -1 0 21690 0 1 64241
box 349 1275 1049 1701
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_6
timestamp 1763476864
transform -1 0 20713 0 1 64241
box 349 1275 1049 1701
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_7
timestamp 1763476864
transform -1 0 42153 0 1 64241
box 349 1275 1049 1701
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_8
timestamp 1763476864
transform -1 0 36525 0 1 64241
box 349 1275 1049 1701
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_9
timestamp 1763476864
transform -1 0 31798 0 1 64241
box 349 1275 1049 1701
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_10
timestamp 1763476864
transform -1 0 40392 0 1 64241
box 349 1275 1049 1701
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_11
timestamp 1763476864
transform -1 0 30900 0 1 64241
box 349 1275 1049 1701
use power_route_512x8m81  power_route_512x8m81_0
timestamp 1763483433
transform 1 0 -1344 0 1 -1785
box 1345 1981 61604 67726
use rcol4_512_512x8m81  rcol4_512_512x8m81_0
timestamp 1763486358
transform 1 0 42157 0 1 3172
box -1076 -2043 17384 62801
use xdec64_512x8m81  xdec64_512x8m81_0
timestamp 1763476864
transform 1 0 20073 0 1 24947
box -2266 -159 21704 39589
<< labels >>
flabel metal3 s 467 22422 467 22422 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 24084 347 24084 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 24947 369 24947 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 25622 347 25622 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 26834 347 26834 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 26159 369 26159 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 27371 369 27371 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 28046 347 28046 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 29258 347 29258 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 28583 369 28583 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 29795 369 29795 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 31007 369 31007 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 32219 369 32219 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 33431 369 33431 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 34643 369 34643 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 35855 369 35855 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 37067 369 37067 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 38279 369 38279 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 45551 369 45551 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 64358 347 64358 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 30422 347 30422 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 31634 347 31634 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 32846 347 32846 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 34058 347 34058 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 35270 347 35270 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 36482 347 36482 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 37694 347 37694 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 63731 369 63731 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 63146 347 63146 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 62519 369 62519 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 61934 347 61934 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 61259 369 61259 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 60722 347 60722 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 60047 369 60047 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 59462 347 59462 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 58835 369 58835 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 58250 347 58250 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 57623 369 57623 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 57038 347 57038 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 56411 369 56411 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 55826 347 55826 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 55199 369 55199 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 54614 347 54614 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 53987 369 53987 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 53402 347 53402 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 52775 369 52775 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 52190 347 52190 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 51563 369 51563 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 50978 347 50978 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 50351 369 50351 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 49766 347 49766 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 48602 347 48602 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 49187 369 49187 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 47390 347 47390 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 47975 369 47975 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 46763 369 46763 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 46178 347 46178 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 44966 347 44966 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 43754 347 43754 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 44339 369 44339 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 42542 347 42542 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 43127 369 43127 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 41330 347 41330 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 41915 369 41915 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 40118 347 40118 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 40703 369 40703 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 39491 369 39491 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 375 38906 375 38906 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 14821 65812 14821 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 18965 65812 18965 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 7893 65812 7893 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 11673 65812 11673 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 7040 65812 7040 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 3260 65812 3260 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 10820 65812 10820 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 65032 369 65032 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 4113 65812 4113 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 21886 65812 21886 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 27399 65812 27399 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 29225 65812 29225 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 25180 65812 25180 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 40672 65812 40672 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 31913 65812 31913 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 32783 65812 32783 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 38373 65812 38373 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 37188 65812 37188 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 34620 65812 34620 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 33637 65812 33637 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 19670 347 19670 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 438 16455 438 16455 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 345 15485 345 15485 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 1375 65812 1375 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 2228 65812 2228 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 13105 65812 13105 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 13958 65812 13958 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 18121 65812 18121 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 17312 65812 17312 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 16451 65812 16451 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 9195 65812 9195 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 10048 65812 10048 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 5285 65812 5285 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 6138 65812 6138 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 21001 65812 21001 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 20024 65812 20024 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 30211 65812 30211 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 31109 65812 31109 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 24327 65812 24327 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 23177 65812 23177 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 26374 65812 26374 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 28427 65812 28427 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 35836 65812 35836 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 39703 65812 39703 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 273 11233 273 11233 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 351 8576 351 8576 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 356 12762 356 12762 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 387 5857 387 5857 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 357 7448 357 7448 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 349 2993 349 2993 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 351 4626 351 4626 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 385 2223 385 2223 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 356 1182 356 1182 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 25571 124 25571 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 27809 124 27809 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 30053 124 30053 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 12839 124 12839 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 6119 124 6119 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 18347 124 18347 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 7799 124 7799 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 13679 124 13679 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 844 124 844 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 22276 124 22276 124 0 FreeSans 313 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 23464 124 23464 124 0 FreeSans 313 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 24732 124 24732 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 26970 124 26970 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 29213 124 29213 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 19257 124 19257 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 1777 124 1777 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 2759 124 2759 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 4439 124 4439 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 5279 124 5279 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 3600 124 3600 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 6958 124 6958 124 0 FreeSans 313 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 11160 124 11160 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 14518 124 14518 124 0 FreeSans 313 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 21077 124 21077 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 9060 124 9060 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 10319 124 10319 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 11999 124 11999 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 20167 124 20167 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 15687 124 15687 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 16527 124 16527 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 17437 124 17437 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 41200 124 41200 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 42110 124 42110 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 39380 124 39380 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 35263 124 35263 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 57062 124 57062 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 34346 124 34346 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 38470 124 38470 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 37085 124 37085 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 31733 124 31733 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 30893 124 30893 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 40290 124 40290 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 32573 124 32573 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 36213 124 36213 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 33413 124 33413 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
rlabel metal2 s 19602 141 19602 141 4 CLK
port 11 nsew signal input
rlabel metal2 s 1380 137 1380 137 4 D[0]
port 19 nsew signal input
rlabel metal2 s 20349 141 20349 141 4 A[8]
port 1 nsew signal input
rlabel metal2 s 20871 141 20871 141 4 A[7]
port 2 nsew signal input
rlabel metal2 s 21679 141 21679 141 4 A[2]
port 7 nsew signal input
rlabel metal2 s 22862 141 22862 141 4 A[1]
port 8 nsew signal input
rlabel metal2 s 24047 141 24047 141 4 A[0]
port 9 nsew signal input
rlabel metal2 s 9970 137 9970 137 4 Q[2]
port 26 nsew signal output
rlabel metal2 s 15694 137 15694 137 4 Q[3]
port 25 nsew signal output
rlabel metal2 s 35318 116 35318 116 4 CEN
port 10 nsew signal input
rlabel metal2 s 38170 147 38170 147 4 A[5]
port 4 nsew signal input
rlabel metal2 s 37720 147 37720 147 4 A[6]
port 3 nsew signal input
rlabel metal2 s 38691 147 38691 147 4 A[4]
port 5 nsew signal input
rlabel metal2 s 16472 137 16472 137 4 WEN[3]
port 35 nsew signal input
rlabel metal2 s 16753 137 16753 137 4 D[3]
port 16 nsew signal input
rlabel metal2 s 8627 137 8627 137 4 D[1]
port 18 nsew signal input
rlabel metal2 s 9499 137 9499 137 4 D[2]
port 17 nsew signal input
rlabel metal2 s 39430 147 39430 147 4 A[3]
port 6 nsew signal input
rlabel metal2 s 8144 137 8144 137 4 Q[1]
port 27 nsew signal output
rlabel metal2 s 9223 137 9223 137 4 WEN[2]
port 36 nsew signal input
rlabel metal2 s 8908 137 8908 137 4 WEN[1]
port 37 nsew signal input
rlabel metal2 s 28508 141 28508 141 4 GWEN
port 20 nsew signal input
rlabel metal2 s 1845 137 1845 137 4 WEN[0]
port 38 nsew signal input
rlabel metal2 s 2484 137 2484 137 4 Q[0]
port 28 nsew signal output
flabel metal3 s 59936 1873 59936 1873 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 60018 22422 60018 22422 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59896 15485 59896 15485 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59988 16455 59988 16455 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59898 19670 59898 19670 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59899 2983 59899 2983 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59902 4616 59902 4616 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59938 5847 59938 5847 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59908 7438 59908 7438 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59902 8566 59902 8566 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59824 11223 59824 11223 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59906 12752 59906 12752 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59906 1182 59906 1182 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59416 124 59416 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 65032 59920 65032 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 43756 124 43756 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 42820 124 42820 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
rlabel metal2 s 43959 137 43959 137 4 Q[4]
port 24 nsew signal output
rlabel metal2 s 43360 137 43360 137 4 WEN[4]
port 34 nsew signal input
rlabel metal2 s 42877 137 42877 137 4 D[4]
port 15 nsew signal input
rlabel metal2 s 50732 137 50732 137 4 WEN[6]
port 32 nsew signal input
rlabel metal2 s 51457 137 51457 137 4 Q[6]
port 22 nsew signal output
rlabel metal2 s 50957 137 50957 137 4 D[6]
port 13 nsew signal input
rlabel metal2 s 50217 137 50217 137 4 WEN[5]
port 33 nsew signal input
rlabel metal2 s 49935 137 49935 137 4 D[5]
port 14 nsew signal input
rlabel metal2 s 49452 137 49452 137 4 Q[5]
port 23 nsew signal output
flabel metal3 s 57843 124 57843 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
rlabel metal2 s 57767 137 57767 137 4 WEN[7]
port 31 nsew signal input
rlabel metal2 s 58223 137 58223 137 4 D[7]
port 12 nsew signal input
rlabel metal2 s 57211 137 57211 137 4 Q[7]
port 21 nsew signal output
flabel metal3 s 52323 65812 52323 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 53177 65812 53177 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 45617 65812 45617 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 49397 65812 49397 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 48543 65812 48543 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 54188 65812 54188 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 44763 65812 44763 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 43321 65812 43321 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 42468 65812 42468 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 47231 65812 47231 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 46378 65812 46378 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 50278 65812 50278 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 51131 65812 51131 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 41464 65812 41464 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 55041 65812 55041 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 56225 65812 56225 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59430 65812 59430 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 58386 65812 58386 65812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 57524 65812 57524 65812 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 52663 124 52663 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 56021 124 56021 124 0 FreeSans 313 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 45942 124 45942 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 46782 124 46782 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 47622 124 47622 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 51822 124 51822 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 53502 124 53502 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 54342 124 54342 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 55182 124 55182 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 45103 124 45103 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 48461 124 48461 124 0 FreeSans 313 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 49102 124 49102 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 50361 124 50361 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59897 63191 59897 63191 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 61979 59897 61979 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 60767 59897 60767 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 59555 59897 59555 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 58343 59897 58343 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 57131 59897 57131 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 55919 59897 55919 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 54707 59897 54707 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 53495 59897 53495 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 52283 59897 52283 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 51071 59897 51071 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 49859 59897 49859 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 48647 59897 48647 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 47435 59897 47435 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 46223 59897 46223 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 45011 59897 45011 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 43799 59897 43799 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 42587 59897 42587 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 41375 59897 41375 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 40163 59897 40163 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 38951 59897 38951 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 37739 59897 37739 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 36527 59897 36527 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 35315 59897 35315 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 34103 59897 34103 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 32891 59897 32891 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 31679 59897 31679 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 30467 59897 30467 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 29255 59897 29255 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 28043 59897 28043 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 26831 59897 26831 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 25619 59897 25619 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59920 57688 59920 57688 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 56476 59920 56476 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 55264 59920 55264 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 54052 59920 54052 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 52840 59920 52840 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 51628 59920 51628 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 50416 59920 50416 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 49204 59920 49204 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 47992 59920 47992 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 46780 59920 46780 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 45568 59920 45568 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 44356 59920 44356 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 43144 59920 43144 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 41932 59920 41932 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 40720 59920 40720 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 39508 59920 39508 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 38296 59920 38296 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 37084 59920 37084 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 35872 59920 35872 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 34660 59920 34660 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 33448 59920 33448 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 32236 59920 32236 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 31024 59920 31024 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 29812 59920 29812 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 28600 59920 28600 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 27388 59920 27388 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 24964 59920 24964 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 26176 59920 26176 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 58900 59920 58900 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 60112 59920 60112 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 61324 59920 61324 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 62536 59920 62536 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 63748 59920 63748 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59897 64383 59897 64383 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 24084 59897 24084 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60260 65973
<< end >>
