magic
tech gf180mcuD
magscale 1 5
timestamp 1763766357
<< metal2 >>
rect -133 14 133 23
rect -133 -14 -125 14
rect 125 -14 133 14
rect -133 -23 133 -14
<< via2 >>
rect -125 -14 125 14
<< metal3 >>
rect -133 14 133 23
rect -133 -14 -125 14
rect 125 -14 133 14
rect -133 -23 133 -14
<< end >>
