magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< nmos >>
rect 0 0 56 318
<< ndiff >>
rect -88 305 0 318
rect -88 13 -75 305
rect -29 13 0 305
rect -88 0 0 13
rect 56 305 144 318
rect 56 13 85 305
rect 131 13 144 305
rect 56 0 144 13
<< ndiffc >>
rect -75 13 -29 305
rect 85 13 131 305
<< polysilicon >>
rect 0 318 56 362
rect 0 -44 56 0
<< metal1 >>
rect -75 305 -29 318
rect -75 0 -29 13
rect 85 305 131 318
rect 85 0 131 13
<< labels >>
flabel ndiffc -40 159 -40 159 0 FreeSans 93 0 0 0 S
flabel ndiffc 96 159 96 159 0 FreeSans 93 0 0 0 D
<< end >>
