magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal2 >>
rect -1299 95 1299 123
rect -1299 -95 -1274 95
rect 1274 -95 1299 95
rect -1299 -122 1299 -95
<< via2 >>
rect -1274 -95 1274 95
<< metal3 >>
rect -1299 95 1299 123
rect -1299 -95 -1274 95
rect 1274 -95 1299 95
rect -1299 -123 1299 -95
<< end >>
