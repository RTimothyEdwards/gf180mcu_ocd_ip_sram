magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< nwell >>
rect -205 0 492 395
<< pmos >>
rect -30 86 318 298
<< pdiff >>
rect -119 277 -30 298
rect -119 231 -105 277
rect -59 231 -30 277
rect -119 153 -30 231
rect -119 107 -105 153
rect -59 107 -30 153
rect -119 86 -30 107
rect 318 277 406 298
rect 318 231 347 277
rect 393 231 406 277
rect 318 153 406 231
rect 318 107 347 153
rect 393 107 406 153
rect 318 86 406 107
<< pdiffc >>
rect -105 231 -59 277
rect -105 107 -59 153
rect 347 231 393 277
rect 347 107 393 153
<< polysilicon >>
rect -30 391 318 404
rect -30 345 -6 391
rect 295 345 318 391
rect -30 298 318 345
rect -30 42 318 86
<< polycontact >>
rect -6 345 295 391
<< metal1 >>
rect -83 391 370 420
rect -83 345 -6 391
rect 295 345 370 391
rect -83 340 370 345
rect -110 277 -56 294
rect -110 231 -105 277
rect -59 231 -56 277
rect -110 153 -56 231
rect -110 107 -105 153
rect -59 107 -56 153
rect -110 25 -56 107
rect 342 277 396 294
rect 342 231 347 277
rect 393 231 396 277
rect 342 153 396 231
rect 342 107 347 153
rect 393 107 396 153
rect 342 25 396 107
rect -127 -131 407 25
rect -110 -132 396 -131
<< end >>
