magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nwell >>
rect -133 -66 160 277
<< polysilicon >>
rect -14 211 41 245
rect -14 -34 41 0
use pmos_5p04310591302014_256x8m81  pmos_5p04310591302014_256x8m81_0
timestamp 1763766357
transform 1 0 -14 0 1 0
box -174 -86 230 297
<< end >>
