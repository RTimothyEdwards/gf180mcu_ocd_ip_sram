magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< polysilicon >>
rect -325 23 325 36
rect -325 -23 -312 23
rect 312 -23 325 23
rect -325 -36 325 -23
<< polycontact >>
rect -312 -23 312 23
<< metal1 >>
rect -319 23 319 30
rect -319 -23 -312 23
rect 312 -23 319 23
rect -319 -30 319 -23
<< end >>
