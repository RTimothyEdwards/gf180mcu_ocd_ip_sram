magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< nwell >>
rect -133 -66 265 489
<< polysilicon >>
rect -42 423 13 456
rect 118 423 173 456
rect -42 -34 13 0
rect 118 -34 173 0
use pmos_5p04310591302058_3v1024x8m81  pmos_5p04310591302058_3v1024x8m81_0
timestamp 1764525316
transform 1 0 -14 0 1 0
box -202 -86 362 509
<< end >>
