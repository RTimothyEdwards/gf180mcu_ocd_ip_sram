magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< nwell >>
rect -154 -530 154 1130
<< nsubdiff >>
rect -53 994 53 1026
rect -53 -394 -23 994
rect 23 -394 53 994
rect -53 -427 53 -394
<< nsubdiffcont >>
rect -23 -394 23 994
<< metal1 >>
rect -40 994 40 1012
rect -40 -394 -23 994
rect 23 -394 40 994
rect -40 -412 40 -394
<< end >>
