magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< error_s >>
rect -201 0 -155 106
rect -41 0 5 106
rect 119 0 165 106
rect 280 0 326 106
rect 440 0 486 106
rect 601 0 647 106
<< polysilicon >>
rect -125 105 -70 140
rect 35 105 90 140
rect 195 105 251 140
rect 356 105 411 140
rect 516 105 572 140
rect -125 -34 -70 0
rect 35 -34 90 0
rect 195 -34 251 0
rect 356 -34 411 0
rect 516 -34 572 0
use nmos_5p04310591302036_512x8m81  nmos_5p04310591302036_512x8m81_0
timestamp 1763476864
transform 1 0 -14 0 1 0
box -200 -44 674 150
<< end >>
