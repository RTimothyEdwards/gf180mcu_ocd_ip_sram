magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< polysilicon >>
rect -95 23 95 36
rect -95 -23 -81 23
rect 81 -23 95 23
rect -95 -36 95 -23
<< polycontact >>
rect -81 -23 81 23
<< metal1 >>
rect -89 23 89 30
rect -89 -23 -81 23
rect 81 -23 89 23
rect -89 -30 89 -23
<< end >>
