magic
tech gf180mcuD
magscale 1 10
timestamp 1763482574
<< metal2 >>
rect 1304 341 1461 481
rect 1777 341 1934 481
rect 2366 341 2522 481
rect 8073 341 8229 481
rect 8544 341 8701 481
rect 8822 341 8979 481
rect 9137 341 9294 481
rect 9417 341 9574 481
rect 9888 341 10045 481
rect 15595 341 15752 481
rect 16382 341 16539 481
rect 16656 341 16813 481
rect 19555 341 19712 481
rect 20304 341 20461 481
rect 20793 341 20950 481
rect 21601 341 21758 481
rect 22786 341 22943 481
rect 23970 341 24126 481
rect 28411 341 28568 481
rect 35239 341 35396 481
rect 37640 341 37797 481
rect 38091 341 38248 481
rect 38614 341 38771 481
rect 39385 341 39542 481
rect 42812 341 42969 481
rect 43280 341 43437 481
rect 43870 341 44027 481
rect 49376 341 49533 481
rect 49847 341 50004 481
rect 50126 341 50282 481
rect 50641 341 50797 481
rect 50921 341 51077 481
rect 51392 341 51548 481
rect 57098 341 57255 481
rect 57686 341 57843 481
rect 58160 341 58317 481
<< metal3 >>
rect 1010 66143 1710 66283
rect 1868 66143 2568 66283
rect 2895 66143 3595 66283
rect 3753 66143 4453 66283
rect 4920 66143 5620 66283
rect 5778 66143 6478 66283
rect 6675 66143 7375 66283
rect 7533 66143 8233 66283
rect 8830 66143 9530 66283
rect 9688 66143 10388 66283
rect 10455 66143 11155 66283
rect 11313 66143 12013 66283
rect 12740 66143 13440 66283
rect 13598 66143 14298 66283
rect 14457 66143 15157 66283
rect 16090 66143 16790 66283
rect 16948 66143 17648 66283
rect 17760 66143 18460 66283
rect 18600 66143 19300 66283
rect 19663 66143 20363 66283
rect 20641 66143 21341 66283
rect 21497 66143 22197 66283
rect 22816 66143 23516 66283
rect 23966 66143 24666 66283
rect 24790 66143 25490 66283
rect 26013 66143 26713 66283
rect 27009 66143 27709 66283
rect 28067 66143 28767 66283
rect 28861 66143 29561 66283
rect 29851 66143 30551 66283
rect 30749 66143 31449 66283
rect 31548 66143 32248 66283
rect 32419 66143 33119 66283
rect 33276 66143 33976 66283
rect 34230 66143 34930 66283
rect 35475 66143 36175 66283
rect 36798 66143 37498 66283
rect 37983 66143 38683 66283
rect 39343 66143 40043 66283
rect 40282 66143 40982 66283
rect 41103 66143 41803 66283
rect 42103 66143 42803 66283
rect 42961 66143 43661 66283
rect 44399 66143 45099 66283
rect 45256 66143 45956 66283
rect 46013 66143 46713 66283
rect 46871 66143 47571 66283
rect 48179 66143 48879 66283
rect 49036 66143 49736 66283
rect 49913 66143 50613 66283
rect 50771 66143 51471 66283
rect 51959 66143 52659 66283
rect 52816 66143 53516 66283
rect 53823 66143 54523 66283
rect 54681 66143 55381 66283
rect 55860 66143 56560 66283
rect 57163 66143 57863 66283
rect 58021 66143 58721 66283
rect 59066 66143 59766 66283
rect 0 65023 140 65723
rect 60120 65024 60260 65723
rect 0 64457 140 64947
rect 60120 64434 60260 64924
rect 0 63827 140 64317
rect 60120 63844 60260 64334
rect 0 63245 140 63735
rect 60120 63242 60260 63732
rect 0 62615 140 63105
rect 60120 62632 60260 63122
rect 0 62033 140 62523
rect 60120 62030 60260 62520
rect 0 61403 140 61893
rect 60120 61420 60260 61910
rect 0 60821 140 61311
rect 60120 60818 60260 61308
rect 0 60191 140 60681
rect 60120 60208 60260 60698
rect 0 59609 140 60099
rect 60120 59606 60260 60096
rect 0 58979 140 59469
rect 60120 58996 60260 59486
rect 0 58397 140 58887
rect 60120 58394 60260 58884
rect 0 57767 140 58257
rect 60120 57784 60260 58274
rect 0 57185 140 57675
rect 60120 57182 60260 57672
rect 0 56555 140 57045
rect 60120 56572 60260 57062
rect 0 55973 140 56463
rect 60120 55970 60260 56460
rect 0 55343 140 55833
rect 60120 55360 60260 55850
rect 0 54761 140 55251
rect 60120 54758 60260 55248
rect 0 54131 140 54621
rect 60120 54148 60260 54638
rect 0 53549 140 54039
rect 60120 53546 60260 54036
rect 0 52919 140 53409
rect 60120 52936 60260 53426
rect 0 52337 140 52827
rect 60120 52334 60260 52824
rect 0 51707 140 52197
rect 60120 51724 60260 52214
rect 0 51125 140 51615
rect 60120 51122 60260 51612
rect 0 50495 140 50985
rect 60120 50512 60260 51002
rect 0 49913 140 50403
rect 60120 49910 60260 50400
rect 0 49283 140 49773
rect 60120 49300 60260 49790
rect 0 48701 140 49191
rect 60120 48698 60260 49188
rect 0 48071 140 48561
rect 60120 48088 60260 48578
rect 0 47489 140 47979
rect 60120 47486 60260 47976
rect 0 46859 140 47349
rect 60120 46876 60260 47366
rect 0 46277 140 46767
rect 60120 46274 60260 46764
rect 0 45647 140 46137
rect 60120 45664 60260 46154
rect 0 45065 140 45555
rect 60120 45062 60260 45552
rect 0 44435 140 44925
rect 60120 44452 60260 44942
rect 0 43853 140 44343
rect 60120 43850 60260 44340
rect 0 43223 140 43713
rect 60120 43240 60260 43730
rect 0 42641 140 43131
rect 60120 42638 60260 43128
rect 0 42011 140 42501
rect 60120 42028 60260 42518
rect 0 41429 140 41919
rect 60120 41426 60260 41916
rect 0 40799 140 41289
rect 60120 40816 60260 41306
rect 0 40217 140 40707
rect 60120 40214 60260 40704
rect 0 39587 140 40077
rect 60120 39604 60260 40094
rect 0 39005 140 39495
rect 60120 39002 60260 39492
rect 0 38375 140 38865
rect 60120 38392 60260 38882
rect 0 37793 140 38283
rect 60120 37790 60260 38280
rect 0 37163 140 37653
rect 60120 37180 60260 37670
rect 0 36581 140 37071
rect 60120 36578 60260 37068
rect 0 35951 140 36441
rect 60120 35968 60260 36458
rect 0 35369 140 35859
rect 60120 35366 60260 35856
rect 0 34739 140 35229
rect 60120 34756 60260 35246
rect 0 34157 140 34647
rect 60120 34154 60260 34644
rect 0 33527 140 34017
rect 60120 33544 60260 34034
rect 0 32945 140 33435
rect 60120 32942 60260 33432
rect 0 32315 140 32805
rect 60120 32332 60260 32822
rect 0 31733 140 32223
rect 60120 31730 60260 32220
rect 0 31103 140 31593
rect 60120 31120 60260 31610
rect 0 30521 140 31011
rect 60120 30518 60260 31008
rect 0 29891 140 30381
rect 60120 29908 60260 30398
rect 0 29309 140 29799
rect 60120 29306 60260 29796
rect 0 28679 140 29169
rect 60120 28696 60260 29186
rect 0 28097 140 28587
rect 60120 28094 60260 28584
rect 0 27467 140 27957
rect 60120 27484 60260 27974
rect 0 26885 140 27375
rect 60120 26882 60260 27372
rect 0 26255 140 26745
rect 60120 26272 60260 26762
rect 0 25673 140 26163
rect 60120 25670 60260 26160
rect 0 25043 140 25533
rect 60120 25060 60260 25550
rect 0 24175 140 24728
rect 60120 24175 60260 24728
rect 0 20940 140 23887
rect 60120 20939 60260 23887
rect 0 19154 140 20541
rect 60120 19154 60260 20541
rect 0 16456 140 17156
rect 60120 16456 60260 17156
rect 0 15297 140 15997
rect 60120 15297 60260 15997
rect 0 12961 140 14867
rect 60120 12951 60260 14857
rect 0 10379 140 12761
rect 60120 10369 60260 12751
rect 0 8775 140 10274
rect 60120 8765 60260 10264
rect 0 7473 140 8395
rect 60120 7463 60260 8385
rect 0 6056 140 7010
rect 60120 6046 60260 7000
rect 0 4386 140 5667
rect 60120 4376 60260 5657
rect 0 3192 140 4290
rect 60120 3182 60260 4280
rect 0 2101 140 2990
rect 60120 2091 60260 2980
rect 0 1203 140 1903
rect 60120 1203 60260 1903
rect 494 341 1194 481
rect 1427 341 2127 481
rect 2409 341 3109 481
rect 3249 341 3949 481
rect 4089 341 4789 481
rect 4929 341 5629 481
rect 5769 341 6469 481
rect 6609 341 7309 481
rect 7449 341 8149 481
rect 8710 341 9410 481
rect 9969 341 10669 481
rect 10809 341 11509 481
rect 11649 341 12349 481
rect 12489 341 13189 481
rect 13329 341 14029 481
rect 14169 341 14869 481
rect 15337 341 16037 481
rect 16177 341 16877 481
rect 17087 341 17787 481
rect 17997 341 18697 481
rect 18907 341 19607 481
rect 19817 341 20517 481
rect 20727 341 21427 481
rect 21926 341 22626 481
rect 23115 341 23815 481
rect 24381 341 25081 481
rect 25221 341 25921 481
rect 26619 341 27319 481
rect 27459 341 28159 481
rect 28863 341 29563 481
rect 29703 341 30403 481
rect 30543 341 31243 481
rect 31383 341 32083 481
rect 32223 341 32923 481
rect 33063 341 33763 481
rect 33996 341 34696 481
rect 34913 341 35613 481
rect 35863 341 36563 481
rect 36734 341 37434 481
rect 38120 341 38820 481
rect 39030 341 39730 481
rect 39940 341 40640 481
rect 40850 341 41550 481
rect 41760 341 42460 481
rect 42670 341 43370 481
rect 43606 341 44306 481
rect 44752 341 45452 481
rect 45592 341 46292 481
rect 46432 341 47132 481
rect 47272 341 47972 481
rect 48112 341 48812 481
rect 48952 341 49652 481
rect 50211 341 50911 481
rect 51472 341 52172 481
rect 52312 341 53012 481
rect 53152 341 53852 481
rect 53992 341 54692 481
rect 54832 341 55532 481
rect 55672 341 56372 481
rect 56712 341 57412 481
rect 57693 341 58393 481
rect 59066 341 59766 481
<< labels >>
flabel metal3 s 70 25963 70 25963 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 25288 70 25288 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 24425 70 24425 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 22763 70 22763 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 26500 70 26500 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 27712 70 27712 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 28924 70 28924 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 30136 70 30136 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 31348 70 31348 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 32560 70 32560 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 33772 70 33772 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 34984 70 34984 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 36196 70 36196 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 37408 70 37408 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 38620 70 38620 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 39832 70 39832 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 41044 70 41044 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 42256 70 42256 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 43468 70 43468 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 44680 70 44680 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 45892 70 45892 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 47104 70 47104 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 48316 70 48316 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 49528 70 49528 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 50740 70 50740 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 51952 70 51952 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 53164 70 53164 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 54376 70 54376 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 55588 70 55588 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 56800 70 56800 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 58012 70 58012 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 59224 70 59224 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 60436 70 60436 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 61648 70 61648 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 62860 70 62860 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 64072 70 64072 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 27127 70 27127 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 28339 70 28339 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 29551 70 29551 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 30763 70 30763 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 31975 70 31975 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 33187 70 33187 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 34399 70 34399 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 35611 70 35611 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 36823 70 36823 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 38035 70 38035 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 39247 70 39247 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 40459 70 40459 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 41671 70 41671 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 42883 70 42883 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 44095 70 44095 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 45307 70 45307 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 46519 70 46519 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 47731 70 47731 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 48943 70 48943 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 50155 70 50155 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 51367 70 51367 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 52579 70 52579 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 53791 70 53791 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 55003 70 55003 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 56215 70 56215 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 57427 70 57427 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 58639 70 58639 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 59851 70 59851 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 61063 70 61063 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 62275 70 62275 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 63487 70 63487 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 64699 70 64699 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 65373 70 65373 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 31898 66218 31898 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 32769 66218 32769 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 40632 66218 40632 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 33626 66218 33626 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 37148 66218 37148 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 38333 66218 38333 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 34580 66218 34580 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 25140 66218 25140 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 7025 66218 7025 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 10805 66218 10805 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 4103 66218 4103 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 11663 66218 11663 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 3245 66218 3245 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 7883 66218 7883 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 27359 66218 27359 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 21847 66218 21847 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 14807 66218 14807 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 18950 66218 18950 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 29211 66218 29211 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 20011 70 20011 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 16796 70 16796 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 15826 70 15826 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 18110 66218 18110 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 16440 66218 16440 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 17298 66218 17298 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 13948 66218 13948 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 13090 66218 13090 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 1360 66218 1360 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 2218 66218 2218 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 10038 66218 10038 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 9180 66218 9180 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 20013 66218 20013 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 20991 66218 20991 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 30201 66218 30201 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 31099 66218 31099 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 28417 66218 28417 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 6128 66218 6128 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 5270 66218 5270 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 23166 66218 23166 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 24316 66218 24316 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 26363 66218 26363 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 35825 66218 35825 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 39693 66218 39693 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 11574 70 11574 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 13103 70 13103 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 8917 70 8917 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 6198 70 6198 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 4967 70 4967 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 3334 70 3334 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 7789 70 7789 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 2564 70 2564 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 1523 70 1523 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 2759 411 2759 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 22276 411 22276 411 0 FreeSans 280 180 0 0 VSS
port 1 nsew
flabel metal3 s 23464 411 23464 411 0 FreeSans 280 180 0 0 VSS
port 1 nsew
flabel metal3 s 24732 411 24732 411 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 26970 411 26970 411 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 29213 411 29213 411 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 844 411 844 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 6958 411 6958 411 0 FreeSans 280 180 0 0 VSS
port 1 nsew
flabel metal3 s 14518 411 14518 411 0 FreeSans 280 180 0 0 VSS
port 1 nsew
flabel metal3 s 20167 411 20167 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 15687 411 15687 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 16527 411 16527 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 17437 411 17437 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 18347 411 18347 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 19257 411 19257 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 1777 411 1777 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 25571 411 25571 411 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 27809 411 27809 411 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 30053 411 30053 411 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 4439 411 4439 411 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 5279 411 5279 411 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 6119 411 6119 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 7799 411 7799 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 9060 411 9060 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 10319 411 10319 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 11999 411 11999 411 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 12839 411 12839 411 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 13679 411 13679 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 3600 411 3600 411 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 21077 411 21077 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 11160 411 11160 411 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 36213 411 36213 411 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 41200 411 41200 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 39380 411 39380 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 40290 411 40290 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 30893 411 30893 411 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 42110 411 42110 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 32573 411 32573 411 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 31733 411 31733 411 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 33413 411 33413 411 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 38470 411 38470 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 34346 411 34346 411 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 37085 411 37085 411 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 35263 411 35263 411 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal2 s 20382 411 20382 411 0 FreeSans 280 0 0 0 A[8]
port 3 nsew
flabel metal2 s 37718 411 37718 411 0 FreeSans 280 0 0 0 A[6]
port 4 nsew
flabel metal2 s 19633 411 19633 411 0 FreeSans 280 0 0 0 CLK
port 5 nsew
flabel metal2 s 1383 411 1383 411 0 FreeSans 280 0 0 0 D[0]
port 6 nsew
flabel metal2 s 20871 411 20871 411 0 FreeSans 280 0 0 0 A[7]
port 7 nsew
flabel metal2 s 21679 411 21679 411 0 FreeSans 280 0 0 0 A[2]
port 8 nsew
flabel metal2 s 22864 411 22864 411 0 FreeSans 280 0 0 0 A[1]
port 9 nsew
flabel metal2 s 24048 411 24048 411 0 FreeSans 280 0 0 0 A[0]
port 10 nsew
flabel metal2 s 9967 411 9967 411 0 FreeSans 280 180 0 0 Q[2]
port 11 nsew
flabel metal2 s 15673 411 15673 411 0 FreeSans 280 180 0 0 Q[3]
port 12 nsew
flabel metal2 s 35317 411 35317 411 0 FreeSans 280 0 0 0 CEN
port 13 nsew
flabel metal2 s 38170 411 38170 411 0 FreeSans 280 0 0 0 A[5]
port 14 nsew
flabel metal2 s 38693 411 38693 411 0 FreeSans 280 0 0 0 A[4]
port 15 nsew
flabel metal2 s 16461 411 16461 411 0 FreeSans 280 180 0 0 WEN[3]
port 16 nsew
flabel metal2 s 16734 411 16734 411 0 FreeSans 280 180 0 0 D[3]
port 19 nsew
flabel metal2 s 8622 411 8622 411 0 FreeSans 280 180 0 0 D[1]
port 20 nsew
flabel metal2 s 9496 411 9496 411 0 FreeSans 280 180 0 0 D[2]
port 21 nsew
flabel metal2 s 39463 411 39463 411 0 FreeSans 280 0 0 0 A[3]
port 22 nsew
flabel metal2 s 8151 411 8151 411 0 FreeSans 280 180 0 0 Q[1]
port 23 nsew
flabel metal2 s 9216 411 9216 411 0 FreeSans 280 180 0 0 WEN[2]
port 28 nsew
flabel metal2 s 8901 411 8901 411 0 FreeSans 280 180 0 0 WEN[1]
port 29 nsew
flabel metal2 s 2444 411 2444 411 0 FreeSans 280 0 0 0 Q[0]
port 36 nsew
flabel metal2 s 28490 411 28490 411 0 FreeSans 280 0 0 0 GWEN
port 37 nsew
flabel metal2 s 1855 411 1855 411 0 FreeSans 280 0 0 0 WEN[0]
port 38 nsew
flabel metal3 s 60196 24425 60196 24425 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 22763 60196 22763 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 65373 60196 65373 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 20011 60196 20011 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 16796 60196 16796 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 15826 60196 15826 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 11564 60196 11564 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 8907 60196 8907 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 4957 60196 4957 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 3730 60196 3730 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 7779 60196 7779 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 6497 60196 6497 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 13093 60196 13093 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 2554 60196 2554 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 1523 60196 1523 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 59416 411 59416 411 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 43756 411 43756 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 57843 411 57843 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 42820 411 42820 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 56862 411 56862 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal2 s 58238 411 58238 411 0 FreeSans 280 180 0 0 D[7]
port 17 nsew
flabel metal2 s 57176 411 57176 411 0 FreeSans 280 180 0 0 Q[7]
port 18 nsew
flabel metal2 s 51470 411 51470 411 0 FreeSans 280 180 0 0 Q[6]
port 24 nsew
flabel metal2 s 43949 411 43949 411 0 FreeSans 280 180 0 0 Q[4]
port 26 nsew
flabel metal2 s 43358 411 43358 411 0 FreeSans 280 180 0 0 WEN[4]
port 30 nsew
flabel metal2 s 57764 411 57764 411 0 FreeSans 280 180 0 0 WEN[7]
port 31 nsew
flabel metal2 s 50719 411 50719 411 0 FreeSans 280 180 0 0 WEN[6]
port 32 nsew
flabel metal2 s 42891 411 42891 411 0 FreeSans 280 180 0 0 D[4]
port 33 nsew
flabel metal2 s 50999 411 50999 411 0 FreeSans 280 180 0 0 D[6]
port 34 nsew
flabel metal2 s 49925 411 49925 411 0 FreeSans 280 180 0 0 D[5]
port 25 nsew
flabel metal2 s 50204 411 50204 411 0 FreeSans 280 180 0 0 WEN[5]
port 27 nsew
flabel metal2 s 49454 411 49454 411 0 FreeSans 280 180 0 0 Q[5]
port 35 nsew
flabel metal3 s 49386 66218 49386 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 53166 66218 53166 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 54173 66218 54173 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 48529 66218 48529 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 52309 66218 52309 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 44749 66218 44749 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 59416 66218 59416 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 45606 66218 45606 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 55031 66218 55031 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 58371 66218 58371 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 57513 66218 57513 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 47221 66218 47221 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 46363 66218 46363 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 43311 66218 43311 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 42453 66218 42453 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 51121 66218 51121 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 50263 66218 50263 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 41453 66218 41453 66218 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 56210 66218 56210 66218 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 55822 411 55822 411 0 FreeSans 280 180 0 0 VSS
port 1 nsew
flabel metal3 s 53302 411 53302 411 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 47422 411 47422 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 49102 411 49102 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 50361 411 50361 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 51622 411 51622 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 46582 411 46582 411 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 45742 411 45742 411 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 54982 411 54982 411 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 54142 411 54142 411 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 48262 411 48262 411 0 FreeSans 280 180 0 0 VSS
port 1 nsew
flabel metal3 s 44902 411 44902 411 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 52462 411 52462 411 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 27172 60196 27172 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 25960 60196 25960 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 28384 60196 28384 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 29596 60196 29596 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 30808 60196 30808 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 32020 60196 32020 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 33232 60196 33232 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 34444 60196 34444 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 35656 60196 35656 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 36868 60196 36868 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 38080 60196 38080 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 39292 60196 39292 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 40504 60196 40504 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 41716 60196 41716 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 42928 60196 42928 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 44140 60196 44140 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 45352 60196 45352 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 46564 60196 46564 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 47776 60196 47776 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 48988 60196 48988 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 50200 60196 50200 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 51412 60196 51412 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 52624 60196 52624 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 53836 60196 53836 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 55048 60196 55048 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 56260 60196 56260 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 57472 60196 57472 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 58684 60196 58684 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 59896 60196 59896 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 61108 60196 61108 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 62320 60196 62320 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 63532 60196 63532 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 61665 60196 61665 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 62877 60196 62877 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 64089 60196 64089 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 64724 60196 64724 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 60453 60196 60453 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 59241 60196 59241 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 58029 60196 58029 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 56817 60196 56817 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 55605 60196 55605 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 54393 60196 54393 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 53181 60196 53181 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 51969 60196 51969 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 50757 60196 50757 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 49545 60196 49545 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 48333 60196 48333 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 47121 60196 47121 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 45909 60196 45909 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 44697 60196 44697 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 43485 60196 43485 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 42273 60196 42273 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 41061 60196 41061 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 39849 60196 39849 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 38637 60196 38637 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 37425 60196 37425 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 36213 60196 36213 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 35001 60196 35001 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 33789 60196 33789 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 32577 60196 32577 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 31365 60196 31365 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 30153 60196 30153 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 28941 60196 28941 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 27729 60196 27729 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 26517 60196 26517 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 25305 60196 25305 0 FreeSans 280 0 0 0 VDD
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 60460 67883
string path 63.580 0.000 63.580 1.000 
<< end >>
