magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< psubdiff >>
rect -29 64519 240 64574
rect -29 64506 239 64519
rect -29 1889 -16 64506
rect 226 1889 239 64506
rect -29 1830 239 1889
<< psubdiffcont >>
rect -16 1889 226 64506
<< metal1 >>
rect -23 64506 233 64513
rect -23 1889 -16 64506
rect 226 1889 233 64506
rect -23 1882 233 1889
<< end >>
