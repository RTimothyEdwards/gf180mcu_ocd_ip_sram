magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -119 324 119 351
rect -119 -324 -93 324
rect 93 -324 119 324
rect -119 -351 119 -324
<< via2 >>
rect -93 -324 93 324
<< metal3 >>
rect -119 324 119 351
rect -119 -324 -93 324
rect 93 -324 119 324
rect -119 -351 119 -324
<< end >>
