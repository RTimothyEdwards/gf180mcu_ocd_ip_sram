magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect -174 -86 230 1737
<< pmos >>
rect 0 0 56 1651
<< pdiff >>
rect -88 1638 0 1651
rect -88 13 -75 1638
rect -29 13 0 1638
rect -88 0 0 13
rect 56 1638 144 1651
rect 56 13 85 1638
rect 131 13 144 1638
rect 56 0 144 13
<< pdiffc >>
rect -75 13 -29 1638
rect 85 13 131 1638
<< polysilicon >>
rect 0 1651 56 1695
rect 0 -44 56 0
<< metal1 >>
rect -75 1638 -29 1651
rect -75 0 -29 13
rect 85 1638 131 1651
rect 85 0 131 13
<< labels >>
flabel pdiffc -40 825 -40 825 0 FreeSans 186 0 0 0 S
flabel pdiffc 96 825 96 825 0 FreeSans 186 0 0 0 D
<< end >>
