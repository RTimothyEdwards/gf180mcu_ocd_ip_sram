magic
tech gf180mcuD
magscale 1 10
timestamp 1765921700
<< metal2 >>
rect -44 562 44 579
rect -44 38 -28 562
rect 28 38 44 562
rect -44 21 44 38
<< via2 >>
rect -28 38 28 562
<< metal3 >>
rect -45 562 45 579
rect -45 38 -28 562
rect 28 38 45 562
rect -45 -119 45 38
<< end >>
