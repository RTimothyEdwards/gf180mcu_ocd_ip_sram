magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect -202 -86 362 245
<< pmos >>
rect -28 0 28 159
rect 132 0 188 159
<< pdiff >>
rect -116 146 -28 159
rect -116 13 -103 146
rect -57 13 -28 146
rect -116 0 -28 13
rect 28 146 132 159
rect 28 13 57 146
rect 103 13 132 146
rect 28 0 132 13
rect 188 146 276 159
rect 188 13 217 146
rect 263 13 276 146
rect 188 0 276 13
<< pdiffc >>
rect -103 13 -57 146
rect 57 13 103 146
rect 217 13 263 146
<< polysilicon >>
rect -28 159 28 203
rect 132 159 188 203
rect -28 -44 28 0
rect 132 -44 188 0
<< metal1 >>
rect -103 146 -57 159
rect -103 0 -57 13
rect 57 146 103 159
rect 57 0 103 13
rect 217 146 263 159
rect 217 0 263 13
<< labels >>
flabel pdiffc 80 79 80 79 0 FreeSans 186 0 0 0 D
flabel pdiffc -68 79 -68 79 0 FreeSans 186 0 0 0 S
flabel pdiffc 228 79 228 79 0 FreeSans 186 0 0 0 S
<< end >>
