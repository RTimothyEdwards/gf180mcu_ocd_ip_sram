magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< psubdiff >>
rect -56 23 56 58
rect -56 -23 -23 23
rect 23 -23 56 23
rect -56 -57 56 -23
<< psubdiffcont >>
rect -23 -23 23 23
<< metal1 >>
rect -49 23 49 51
rect -49 -23 -23 23
rect 23 -23 49 23
rect -49 -51 49 -23
<< end >>
