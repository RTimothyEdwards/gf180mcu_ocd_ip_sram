magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -119 172 119 198
rect -119 -172 -93 172
rect 93 -172 119 172
rect -119 -198 119 -172
<< via2 >>
rect -93 -172 93 172
<< metal3 >>
rect -119 172 119 198
rect -119 -172 -93 172
rect 93 -172 119 172
rect -119 -198 119 -172
<< end >>
