magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nmos >>
rect -28 0 28 308
rect 132 0 188 308
<< ndiff >>
rect -116 295 -28 308
rect -116 13 -103 295
rect -57 13 -28 295
rect -116 0 -28 13
rect 28 295 132 308
rect 28 13 57 295
rect 103 13 132 295
rect 28 0 132 13
rect 188 295 276 308
rect 188 13 217 295
rect 263 13 276 295
rect 188 0 276 13
<< ndiffc >>
rect -103 13 -57 295
rect 57 13 103 295
rect 217 13 263 295
<< polysilicon >>
rect -28 308 28 352
rect 132 308 188 352
rect -28 -44 28 0
rect 132 -44 188 0
<< metal1 >>
rect -103 295 -57 308
rect -103 0 -57 13
rect 57 295 103 308
rect 57 0 103 13
rect 217 295 263 308
rect 217 0 263 13
<< labels >>
flabel ndiffc 80 154 80 154 0 FreeSans 93 0 0 0 D
flabel ndiffc -68 154 -68 154 0 FreeSans 93 0 0 0 S
flabel ndiffc 227 154 227 154 0 FreeSans 93 0 0 0 S
<< end >>
