magic
tech gf180mcuD
magscale 1 10
timestamp 1763575302
<< metal2 >>
rect -113 467 113 474
rect -113 -627 -106 467
rect 106 -627 113 467
rect -113 -634 113 -627
<< via2 >>
rect -106 -627 106 467
<< metal3 >>
rect -113 467 113 474
rect -113 -627 -106 467
rect 106 -627 113 467
rect -113 -634 113 -627
<< end >>
