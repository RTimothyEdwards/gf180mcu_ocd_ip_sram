magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< nwell >>
rect -18 611 5184 2069
<< pdiff >>
rect 1287 710 1350 844
rect 1548 710 1634 844
rect 3054 710 3104 1030
rect 3299 896 3324 1030
<< polysilicon >>
rect 1409 2288 1465 2374
rect 1569 2288 1625 2374
rect 181 1582 237 2209
rect 341 1582 397 2209
rect 502 1582 558 2209
rect 1409 2102 1465 2211
rect 1569 2102 1625 2211
rect 1730 2102 1786 2219
rect 1890 2102 1946 2219
rect 2051 2102 2107 2219
rect 2211 2102 2267 2219
rect 2372 2102 2428 2219
rect 2532 2102 2588 2219
rect 2693 2102 2749 2219
rect 2853 2102 2909 2219
rect 1124 2044 2909 2102
rect 1124 1969 1249 2044
rect 1409 1874 1465 2044
rect 1569 1874 1625 2044
rect 1730 1874 1786 2044
rect 1890 1874 1946 2044
rect 2051 1874 2107 2044
rect 2211 1874 2267 2044
rect 2372 1874 2428 2044
rect 2532 1874 2588 2044
rect 2693 1874 2749 2044
rect 2853 1874 2909 2044
rect 3270 1878 3326 2213
rect 3430 1878 3486 2213
rect 3591 1878 3647 2213
rect 3751 1878 3807 2213
rect 3912 1878 3968 2213
rect 4072 1878 4128 2213
rect 4233 1878 4289 2213
rect 4393 1878 4449 2213
rect 4554 1878 4610 2213
rect 4714 1878 4770 2213
rect 181 1293 237 1362
rect 341 1293 397 1362
rect 502 1293 558 1362
rect 662 1293 718 1362
rect 823 1293 879 1362
rect 983 1293 1039 1362
rect 3270 1316 3326 1354
rect 3430 1316 3486 1354
rect 3591 1316 3647 1354
rect 3751 1316 3807 1354
rect 3912 1316 3968 1354
rect 4072 1316 4128 1354
rect 4233 1316 4289 1354
rect 4393 1316 4449 1354
rect 4554 1316 4610 1354
rect 4714 1316 4770 1354
rect 176 1234 1044 1293
rect 3270 1266 4770 1316
rect 3270 1249 4767 1266
rect 1417 1184 1473 1185
rect 846 1141 1473 1184
rect 366 965 422 1077
rect 846 962 902 1141
rect 1417 842 1473 1141
rect 2777 1075 2993 1133
rect 2777 962 2833 1075
rect 2937 962 2993 1075
rect 3157 1068 3213 1175
rect 3411 1068 3467 1249
rect 366 400 422 673
rect 526 400 582 673
rect 846 630 902 671
rect 830 558 902 630
rect 961 625 1361 668
rect 846 455 902 558
rect 1298 599 1361 625
rect 1672 653 1728 671
rect 1298 556 1568 599
rect 1512 508 1568 556
rect 1672 581 1748 653
rect 1672 508 1728 581
rect 1983 509 2037 670
rect 2317 498 2373 673
rect 2477 498 2533 673
rect 3411 620 3467 778
rect 3728 638 3784 667
rect 3888 638 3944 667
rect 4049 638 4105 667
rect 4209 638 4265 667
rect 4370 638 4426 667
rect 4530 638 4586 667
rect 4692 638 4748 667
rect 3728 635 4748 638
rect 3392 571 3467 620
rect 3727 586 4748 635
rect 3392 470 3448 571
rect 3727 511 3783 586
rect 3887 511 3943 586
rect 4048 511 4104 586
rect 4208 511 4264 586
rect 4369 511 4425 586
rect 4529 511 4585 586
rect 4690 511 4746 586
rect 526 196 582 229
rect 846 142 902 283
rect 1983 222 2039 339
rect 1707 163 2039 222
rect 2317 222 2373 305
rect 2477 222 2533 307
rect 2317 163 2533 222
rect 1154 142 1210 160
rect 846 69 1210 142
rect 2777 125 2833 155
rect 2937 125 2993 155
rect 3232 144 3288 296
rect 2777 80 2993 125
rect 2777 79 2833 80
rect 1154 -61 1210 69
<< metal1 >>
rect 265 2016 313 2362
rect 586 2016 634 2354
rect 1499 2142 1545 2420
rect 1819 2142 1866 2364
rect 2141 2142 2188 2363
rect 2460 2142 2507 2363
rect 2783 2142 2830 2352
rect 977 2093 2830 2142
rect 265 1969 1214 2016
rect 265 1532 313 1969
rect 586 1536 634 1969
rect 907 1543 956 1969
rect 1499 1582 1545 2093
rect 1819 1583 1866 2093
rect 1834 1582 1866 1583
rect 2141 1582 2188 2093
rect 2460 1582 2507 2093
rect 2783 1582 2830 2093
rect 3351 2134 3398 2356
rect 3672 2134 3721 2354
rect 3991 2134 4039 2358
rect 4313 2134 4362 2357
rect 4633 2134 4681 2356
rect 3351 2085 4681 2134
rect 3351 1582 3398 2085
rect 3672 1582 3721 2085
rect 3991 1582 4039 2085
rect 4313 1582 4362 2085
rect 4633 1582 4681 2085
rect 321 1085 434 1267
rect 611 1225 3045 1274
rect 611 908 657 1225
rect 2401 1178 2450 1179
rect 930 1138 962 1142
rect 930 1111 979 1138
rect 290 16 339 755
rect 610 624 658 751
rect 744 716 835 1022
rect 610 565 773 624
rect 610 269 658 565
rect 931 116 979 1111
rect 2401 1131 2909 1178
rect 1100 267 1190 1022
rect 1257 844 1346 1022
rect 1596 845 1643 1022
rect 1257 710 1403 844
rect 1533 710 1643 845
rect 1736 716 1826 1022
rect 1257 507 1346 710
rect 1257 386 1508 507
rect 1596 387 1643 710
rect 1913 641 1964 1022
rect 2050 716 2139 1022
rect 1806 593 1964 641
rect 1609 386 1641 387
rect 1257 216 1346 386
rect 1913 216 1964 593
rect 2401 387 2450 1131
rect 2683 654 2772 1022
rect 2859 970 2909 1131
rect 2996 1094 3045 1225
rect 2869 716 2901 970
rect 3026 893 3132 1027
rect 3261 893 3398 1028
rect 3026 654 3086 893
rect 3465 716 3554 1022
rect 3633 716 3723 1022
rect 2683 640 3086 654
rect 3792 654 3873 1263
rect 3946 716 4036 1022
rect 4106 654 4186 1260
rect 4260 716 4350 1022
rect 4419 654 4500 1260
rect 4573 716 4664 1022
rect 4733 655 4792 1263
rect 4733 654 4813 655
rect 3157 640 3203 641
rect 2683 586 3692 640
rect 2683 570 3086 586
rect 1257 169 1826 216
rect 1913 169 2424 216
rect 2683 201 2772 570
rect 2839 201 2929 507
rect 2996 201 3086 570
rect 3157 396 3203 586
rect 3792 570 4813 654
rect 3792 392 3873 570
rect 4106 392 4186 570
rect 4419 392 4500 570
rect 4760 386 4813 570
rect 931 69 2884 116
rect 3229 -4 3275 146
rect 1211 -52 3275 -4
<< metal2 >>
rect 1100 266 1190 1022
rect 1101 35 1190 266
rect 2839 201 2929 1022
rect 3308 201 3397 1022
rect 261 -6 1190 35
rect 261 -21 1188 -6
<< metal3 >>
rect 63 2289 5184 2488
rect 1402 1924 1674 1985
rect 63 1396 5184 1595
rect 883 1111 3339 1173
rect 63 710 5184 1028
rect 63 262 5184 507
rect 513 94 603 186
use M1_NACTIVE4310591302028_512x8m81  M1_NACTIVE4310591302028_512x8m81_0
timestamp 1763765945
transform 1 0 1223 0 1 1492
box -36 -95 36 95
use M1_NACTIVE4310591302028_512x8m81  M1_NACTIVE4310591302028_512x8m81_1
timestamp 1763765945
transform 1 0 3089 0 1 1492
box -36 -95 36 95
use M1_NACTIVE4310591302070_512x8m81  M1_NACTIVE4310591302070_512x8m81_0
timestamp 1763765945
transform 1 0 4984 0 1 1492
box -62 -95 62 95
use M1_NACTIVE_01_512x8m81  M1_NACTIVE_01_512x8m81_0
timestamp 1763765945
transform 1 0 4986 0 1 876
box -53 -112 53 113
use M1_NACTIVE_01_512x8m81  M1_NACTIVE_01_512x8m81_2
timestamp 1763765945
transform 1 0 109 0 1 876
box -53 -112 53 113
use M1_PACTIVE4310591302039_512x8m81  M1_PACTIVE4310591302039_512x8m81_0
timestamp 1763765945
transform 1 0 3089 0 1 2385
box -36 -95 36 95
use M1_PACTIVE4310591302069_512x8m81  M1_PACTIVE4310591302069_512x8m81_0
timestamp 1763765945
transform 1 0 4984 0 1 381
box -62 -95 62 95
use M1_PACTIVE4310591302069_512x8m81  M1_PACTIVE4310591302069_512x8m81_1
timestamp 1763765945
transform 1 0 4984 0 1 2385
box -62 -95 62 95
use M1_PACTIVE4310591302071_512x8m81  M1_PACTIVE4310591302071_512x8m81_0
timestamp 1763765945
transform 1 0 998 0 1 2385
box -128 -95 128 95
use M1_PACTIVE_01_512x8m81  M1_PACTIVE_01_512x8m81_0
timestamp 1763765945
transform 1 0 109 0 1 385
box -53 -112 53 113
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_0
timestamp 1763765945
transform 1 0 2827 0 1 92
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_1
timestamp 1763765945
transform 1 0 3035 0 1 1107
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_2
timestamp 1763765945
transform 1 0 3670 0 1 616
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_3
timestamp 1763765945
transform 1 0 3833 0 1 1239
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_4
timestamp 1763765945
transform 1 0 3254 0 1 148
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_5
timestamp 1763765945
transform 1 0 3274 0 1 1139
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_6
timestamp 1763765945
transform 1 0 4143 0 1 1239
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_7
timestamp 1763765945
transform 1 0 4461 0 1 1239
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_8
timestamp 1763765945
transform 1 0 4701 0 1 1239
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_9
timestamp 1763765945
transform 0 -1 988 1 0 605
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_10
timestamp 1763765945
transform 1 0 575 0 1 162
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_11
timestamp 1763765945
transform 1 0 770 0 1 594
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_12
timestamp 1763765945
transform 1 0 1805 0 1 617
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_13
timestamp 1763765945
transform 1 0 1769 0 1 192
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_14
timestamp 1763765945
transform 1 0 2367 0 1 192
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_15
timestamp 1763765945
transform 1 0 1243 0 1 -26
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_16
timestamp 1763765945
transform 1 0 378 0 1 1244
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_17
timestamp 1763765945
transform 1 0 378 0 1 1104
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_18
timestamp 1763765945
transform 1 0 1187 0 1 1992
box -62 -36 62 36
use M2_M1$$201262124_512x8m81  M2_M1$$201262124_512x8m81_0
timestamp 1763765945
transform 1 0 561 0 1 140
box -119 -46 119 46
use M2_M1$$202395692_512x8m81  M2_M1$$202395692_512x8m81_0
timestamp 1763765945
transform 1 0 3509 0 1 395
box -44 -111 44 112
use M2_M1$$202395692_512x8m81  M2_M1$$202395692_512x8m81_1
timestamp 1763765945
transform 1 0 790 0 1 395
box -44 -111 44 112
use M2_M1$$202395692_512x8m81  M2_M1$$202395692_512x8m81_2
timestamp 1763765945
transform 1 0 1781 0 1 395
box -44 -111 44 112
use M2_M1$$202395692_512x8m81  M2_M1$$202395692_512x8m81_3
timestamp 1763765945
transform 1 0 2095 0 1 395
box -44 -111 44 112
use M2_M1$$202396716_512x8m81  M2_M1$$202396716_512x8m81_0
timestamp 1763765945
transform 1 0 1145 0 1 612
box -44 -351 44 351
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_0
timestamp 1763765945
transform 1 0 3678 0 -1 875
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_1
timestamp 1763765945
transform 1 0 2884 0 1 869
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_2
timestamp 1763765945
transform 1 0 4986 0 1 876
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_3
timestamp 1763765945
transform 1 0 4619 0 1 385
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_4
timestamp 1763765945
transform 1 0 4305 0 1 385
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_5
timestamp 1763765945
transform 1 0 3992 0 1 385
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_6
timestamp 1763765945
transform 1 0 3678 0 1 385
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_7
timestamp 1763765945
transform 1 0 3509 0 1 869
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_8
timestamp 1763765945
transform 1 0 3353 0 1 355
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_9
timestamp 1763765945
transform 1 0 3353 0 1 869
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_10
timestamp 1763765945
transform 1 0 2884 0 1 355
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_11
timestamp 1763765945
transform 1 0 3992 0 -1 875
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_12
timestamp 1763765945
transform 1 0 4305 0 -1 875
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_13
timestamp 1763765945
transform 1 0 4619 0 -1 875
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_14
timestamp 1763765945
transform 1 0 1781 0 1 869
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_15
timestamp 1763765945
transform 1 0 2095 0 1 869
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_16
timestamp 1763765945
transform 1 0 109 0 1 876
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_17
timestamp 1763765945
transform 1 0 109 0 1 385
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_18
timestamp 1763765945
transform 1 0 476 0 1 869
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_19
timestamp 1763765945
transform 1 0 476 0 1 385
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_20
timestamp 1763765945
transform 1 0 790 0 1 869
box -45 -122 45 123
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_0
timestamp 1763765945
transform 0 -1 3276 1 0 1142
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_1
timestamp 1763765945
transform 0 -1 319 1 0 14
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_2
timestamp 1763765945
transform 0 -1 946 1 0 1142
box -34 -63 34 63
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_0
timestamp 1763765945
transform 1 0 2582 0 1 882
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_1
timestamp 1763765945
transform 1 0 2582 0 1 372
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_2
timestamp 1763765945
transform 1 0 2268 0 1 882
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_3
timestamp 1763765945
transform 1 0 2268 0 1 372
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_4
timestamp 1763765945
transform 1 0 2320 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_5
timestamp 1763765945
transform 1 0 1379 0 1 2389
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_6
timestamp 1763765945
transform 1 0 1693 0 1 2389
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_7
timestamp 1763765945
transform 1 0 2006 0 1 2389
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_8
timestamp 1763765945
transform 1 0 2320 0 1 2389
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_9
timestamp 1763765945
transform 1 0 1223 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_10
timestamp 1763765945
transform 1 0 140 0 1 2389
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_11
timestamp 1763765945
transform 1 0 453 0 1 2389
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_12
timestamp 1763765945
transform 1 0 453 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_13
timestamp 1763765945
transform 1 0 140 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_14
timestamp 1763765945
transform 1 0 1080 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_15
timestamp 1763765945
transform 1 0 767 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_16
timestamp 1763765945
transform 1 0 2006 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_17
timestamp 1763765945
transform 1 0 1693 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_18
timestamp 1763765945
transform 1 0 1379 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_19
timestamp 1763765945
transform 1 0 4486 0 1 2389
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_20
timestamp 1763765945
transform 1 0 3089 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_21
timestamp 1763765945
transform 1 0 3089 0 1 2389
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_22
timestamp 1763765945
transform 1 0 2947 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_23
timestamp 1763765945
transform 1 0 2634 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_24
timestamp 1763765945
transform 1 0 2947 0 1 2389
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_25
timestamp 1763765945
transform 1 0 2634 0 1 2389
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_26
timestamp 1763765945
transform 1 0 3859 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_27
timestamp 1763765945
transform 1 0 3545 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_28
timestamp 1763765945
transform 1 0 3231 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_29
timestamp 1763765945
transform 1 0 4172 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_30
timestamp 1763765945
transform 1 0 4799 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_31
timestamp 1763765945
transform 1 0 4486 0 1 1495
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_32
timestamp 1763765945
transform 1 0 3231 0 1 2389
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_33
timestamp 1763765945
transform 1 0 3545 0 1 2389
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_34
timestamp 1763765945
transform 1 0 3859 0 1 2389
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_35
timestamp 1763765945
transform 1 0 4172 0 1 2389
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_36
timestamp 1763765945
transform 1 0 4799 0 1 2389
box -34 -99 34 99
use M2_M14310591302025_512x8m81  M2_M14310591302025_512x8m81_0
timestamp 1763765945
transform 0 -1 1538 1 0 1959
box -34 -85 34 135
use M2_M14310591302073_512x8m81  M2_M14310591302073_512x8m81_0
timestamp 1763765945
transform 1 0 4989 0 1 384
box -63 -99 63 99
use M2_M14310591302073_512x8m81  M2_M14310591302073_512x8m81_1
timestamp 1763765945
transform 1 0 4989 0 1 2389
box -63 -99 63 99
use M2_M14310591302073_512x8m81  M2_M14310591302073_512x8m81_2
timestamp 1763765945
transform 1 0 4985 0 1 1495
box -63 -99 63 99
use M2_M14310591302074_512x8m81  M2_M14310591302074_512x8m81_0
timestamp 1763765945
transform 1 0 1003 0 1 2389
box -99 -99 99 99
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_0
timestamp 1763765945
transform 1 0 3678 0 -1 875
box -45 -122 45 123
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_1
timestamp 1763765945
transform 1 0 4619 0 1 385
box -45 -122 45 123
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_2
timestamp 1763765945
transform 1 0 4986 0 1 876
box -45 -122 45 123
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_3
timestamp 1763765945
transform 1 0 3678 0 1 385
box -45 -122 45 123
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_4
timestamp 1763765945
transform 1 0 3992 0 1 385
box -45 -122 45 123
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_5
timestamp 1763765945
transform 1 0 4305 0 1 385
box -45 -122 45 123
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_6
timestamp 1763765945
transform 1 0 3509 0 1 869
box -45 -122 45 123
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_7
timestamp 1763765945
transform 1 0 3992 0 -1 875
box -45 -122 45 123
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_8
timestamp 1763765945
transform 1 0 4619 0 -1 875
box -45 -122 45 123
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_9
timestamp 1763765945
transform 1 0 4305 0 -1 875
box -45 -122 45 123
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_10
timestamp 1763765945
transform 1 0 1781 0 1 869
box -45 -122 45 123
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_11
timestamp 1763765945
transform 1 0 2095 0 1 869
box -45 -122 45 123
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_12
timestamp 1763765945
transform 1 0 109 0 1 876
box -45 -122 45 123
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_13
timestamp 1763765945
transform 1 0 109 0 1 385
box -45 -122 45 123
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_14
timestamp 1763765945
transform 1 0 476 0 1 869
box -45 -122 45 123
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_15
timestamp 1763765945
transform 1 0 476 0 1 385
box -45 -122 45 123
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_16
timestamp 1763765945
transform 1 0 790 0 1 869
box -45 -122 45 123
use M3_M2$$201255980_512x8m81  M3_M2$$201255980_512x8m81_0
timestamp 1763765945
transform 1 0 561 0 1 139
box -119 -46 119 46
use M3_M2$$202397740_512x8m81  M3_M2$$202397740_512x8m81_0
timestamp 1763765945
transform 1 0 3509 0 1 395
box -45 -112 45 112
use M3_M2$$202397740_512x8m81  M3_M2$$202397740_512x8m81_1
timestamp 1763765945
transform 1 0 1781 0 1 395
box -45 -112 45 112
use M3_M2$$202397740_512x8m81  M3_M2$$202397740_512x8m81_2
timestamp 1763765945
transform 1 0 2095 0 1 395
box -45 -112 45 112
use M3_M2$$202397740_512x8m81  M3_M2$$202397740_512x8m81_3
timestamp 1763765945
transform 1 0 790 0 1 385
box -45 -112 45 112
use M3_M2431059130207_512x8m81  M3_M2431059130207_512x8m81_0
timestamp 1763765945
transform 1 0 3276 0 1 1142
box -63 -35 63 35
use M3_M2431059130207_512x8m81  M3_M2431059130207_512x8m81_1
timestamp 1763765945
transform 1 0 946 0 1 1142
box -63 -35 63 35
use M3_M24310591302026_512x8m81  M3_M24310591302026_512x8m81_0
timestamp 1763765945
transform 0 -1 1538 1 0 1959
box -35 -135 35 135
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_0
timestamp 1763765945
transform 1 0 2582 0 1 882
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_1
timestamp 1763765945
transform 1 0 2582 0 1 372
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_2
timestamp 1763765945
transform 1 0 2268 0 1 882
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_3
timestamp 1763765945
transform 1 0 2268 0 1 372
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_4
timestamp 1763765945
transform 1 0 1080 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_5
timestamp 1763765945
transform 1 0 767 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_6
timestamp 1763765945
transform 1 0 1223 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_7
timestamp 1763765945
transform 1 0 453 0 1 2389
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_8
timestamp 1763765945
transform 1 0 1379 0 1 2389
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_9
timestamp 1763765945
transform 1 0 1693 0 1 2389
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_10
timestamp 1763765945
transform 1 0 2006 0 1 2389
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_11
timestamp 1763765945
transform 1 0 2320 0 1 2389
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_12
timestamp 1763765945
transform 1 0 140 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_13
timestamp 1763765945
transform 1 0 140 0 1 2389
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_14
timestamp 1763765945
transform 1 0 453 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_15
timestamp 1763765945
transform 1 0 1379 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_16
timestamp 1763765945
transform 1 0 1693 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_17
timestamp 1763765945
transform 1 0 2006 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_18
timestamp 1763765945
transform 1 0 2320 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_19
timestamp 1763765945
transform 1 0 2947 0 1 2389
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_20
timestamp 1763765945
transform 1 0 2634 0 1 2389
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_21
timestamp 1763765945
transform 1 0 3231 0 1 2389
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_22
timestamp 1763765945
transform 1 0 3545 0 1 2389
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_23
timestamp 1763765945
transform 1 0 3859 0 1 2389
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_24
timestamp 1763765945
transform 1 0 4172 0 1 2389
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_25
timestamp 1763765945
transform 1 0 4799 0 1 2389
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_26
timestamp 1763765945
transform 1 0 4486 0 1 2389
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_27
timestamp 1763765945
transform 1 0 2947 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_28
timestamp 1763765945
transform 1 0 2634 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_29
timestamp 1763765945
transform 1 0 3231 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_30
timestamp 1763765945
transform 1 0 3545 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_31
timestamp 1763765945
transform 1 0 3859 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_32
timestamp 1763765945
transform 1 0 4172 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_33
timestamp 1763765945
transform 1 0 4799 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_34
timestamp 1763765945
transform 1 0 4486 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_35
timestamp 1763765945
transform 1 0 3089 0 1 1495
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_36
timestamp 1763765945
transform 1 0 3089 0 1 2389
box -35 -99 35 99
use M3_M24310591302050_512x8m81  M3_M24310591302050_512x8m81_0
timestamp 1763765945
transform 1 0 1003 0 1 2389
box -99 -99 99 99
use M3_M24310591302072_512x8m81  M3_M24310591302072_512x8m81_0
timestamp 1763765945
transform 1 0 4989 0 1 384
box -63 -99 63 99
use M3_M24310591302072_512x8m81  M3_M24310591302072_512x8m81_1
timestamp 1763765945
transform 1 0 4989 0 1 2389
box -63 -99 63 99
use M3_M24310591302072_512x8m81  M3_M24310591302072_512x8m81_2
timestamp 1763765945
transform 1 0 4985 0 1 1495
box -63 -99 63 99
use nmos_1p2$$202595372_512x8m81  nmos_1p2$$202595372_512x8m81_0
timestamp 1763765945
transform 1 0 1997 0 1 380
box -102 -44 130 133
use nmos_1p2$$202595372_512x8m81  nmos_1p2$$202595372_512x8m81_1
timestamp 1763765945
transform 1 0 1526 0 1 380
box -102 -44 130 133
use nmos_1p2$$202596396_512x8m81  nmos_1p2$$202596396_512x8m81_0
timestamp 1763765945
transform 1 0 1686 0 1 380
box -102 -44 130 133
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_0
timestamp 1763765945
transform 1 0 3392 0 -1 428
box -88 -44 144 133
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_1
timestamp 1763765945
transform 1 0 3232 0 -1 428
box -88 -44 144 133
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_2
timestamp 1763765945
transform 1 0 366 0 1 269
box -88 -44 144 133
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_3
timestamp 1763765945
transform 1 0 526 0 1 269
box -88 -44 144 133
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_4
timestamp 1763765945
transform 1 0 846 0 1 326
box -88 -44 144 133
use nmos_5p04310591302010_512x8m81  nmos_5p04310591302010_512x8m81_0
timestamp 1763765945
transform 1 0 1154 0 1 196
box -88 -44 144 255
use nmos_5p04310591302039_512x8m81  nmos_5p04310591302039_512x8m81_0
timestamp 1763765945
transform 1 0 2805 0 1 196
box -116 -44 276 255
use nmos_5p04310591302075_512x8m81  nmos_5p04310591302075_512x8m81_0
timestamp 1763765945
transform 1 0 3522 0 1 2249
box -340 -44 1336 223
use nmos_5p04310591302075_512x8m81  nmos_5p04310591302075_512x8m81_1
timestamp 1763765945
transform 1 0 1661 0 1 2249
box -340 -44 1336 223
use nmos_5p04310591302076_512x8m81  nmos_5p04310591302076_512x8m81_0
timestamp 1763765945
transform 1 0 2345 0 1 346
box -116 -44 276 156
use nmos_5p04310591302078_512x8m81  nmos_5p04310591302078_512x8m81_0
timestamp 1763765945
transform 1 0 285 0 1 2249
box -192 -44 361 230
use nmos_5p04310591302081_512x8m81  nmos_5p04310591302081_512x8m81_0
timestamp 1763765945
transform 1 0 3895 0 1 386
box -256 -44 939 128
use pmos_1p2$$202586156_512x8m81  pmos_1p2$$202586156_512x8m81_0
timestamp 1763765945
transform 1 0 1686 0 1 710
box -188 -86 216 297
use pmos_1p2$$202587180_512x8m81  pmos_1p2$$202587180_512x8m81_0
timestamp 1763765945
transform 1 0 1176 0 1 710
box -188 -86 216 297
use pmos_5p04310591302014_512x8m81  pmos_5p04310591302014_512x8m81_0
timestamp 1763765945
transform 1 0 3411 0 -1 1030
box -174 -86 230 297
use pmos_5p04310591302014_512x8m81  pmos_5p04310591302014_512x8m81_1
timestamp 1763765945
transform 1 0 526 0 1 710
box -174 -86 230 297
use pmos_5p04310591302014_512x8m81  pmos_5p04310591302014_512x8m81_2
timestamp 1763765945
transform 1 0 1982 0 1 710
box -174 -86 230 297
use pmos_5p04310591302014_512x8m81  pmos_5p04310591302014_512x8m81_3
timestamp 1763765945
transform 1 0 366 0 1 710
box -174 -86 230 297
use pmos_5p04310591302014_512x8m81  pmos_5p04310591302014_512x8m81_4
timestamp 1763765945
transform 1 0 846 0 1 710
box -174 -86 230 297
use pmos_5p04310591302020_512x8m81  pmos_5p04310591302020_512x8m81_0
timestamp 1763765945
transform 1 0 2805 0 1 710
box -202 -86 362 297
use pmos_5p04310591302041_512x8m81  pmos_5p04310591302041_512x8m81_0
timestamp 1763765945
transform 1 0 3157 0 -1 1030
box -174 -86 230 175
use pmos_5p04310591302041_512x8m81  pmos_5p04310591302041_512x8m81_1
timestamp 1763765945
transform 1 0 1417 0 1 710
box -174 -86 230 175
use pmos_5p04310591302077_512x8m81  pmos_5p04310591302077_512x8m81_0
timestamp 1763765945
transform 1 0 1661 0 1 1398
box -426 -86 1422 526
use pmos_5p04310591302077_512x8m81  pmos_5p04310591302077_512x8m81_2
timestamp 1763765945
transform 1 0 3522 0 1 1398
box -426 -86 1422 526
use pmos_5p04310591302079_512x8m81  pmos_5p04310591302079_512x8m81_0
timestamp 1763765945
transform 1 0 3884 0 1 710
box -330 -86 1038 291
use pmos_5p04310591302080_512x8m81  pmos_5p04310591302080_512x8m81_0
timestamp 1763765945
transform 1 0 2345 0 1 710
box -202 -86 362 351
use pmos_5p04310591302082_512x8m81  pmos_5p04310591302082_512x8m81_0
timestamp 1763765945
transform 1 0 321 0 1 1398
box -314 -86 892 317
<< labels >>
rlabel metal3 s 176 2435 176 2435 4 vss
port 1 nsew
rlabel metal3 s 176 1522 176 1522 4 vdd
port 3 nsew
rlabel metal1 s 4644 2102 4644 2102 4 GWE
port 6 nsew
rlabel metal1 s 336 1119 336 1119 4 wen
port 5 nsew
rlabel metal3 s 605 162 605 162 4 clk
port 4 nsew
rlabel metal3 s 176 869 176 869 4 vdd
port 3 nsew
rlabel metal3 s 176 385 176 385 4 vss
port 1 nsew
flabel metal3 s 1537 1955 1537 1955 0 FreeSans 700 0 0 0 IGWEN
port 2 nsew
<< properties >>
string path 6.310 7.305 23.850 7.305 
<< end >>
