magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< error_s >>
rect 439 5562 440 5948
rect 255 5506 294 5562
rect 384 5506 440 5562
rect 311 5488 350 5506
rect 384 5488 423 5506
rect 439 5488 440 5506
rect 456 5488 495 5506
rect 529 5488 568 5562
rect 764 5510 803 5566
rect 820 5492 859 5510
rect 893 5492 932 5566
<< nwell >>
rect 300 1924 389 2148
<< polysilicon >>
rect 525 5252 580 5279
rect 525 5240 589 5252
rect 533 5153 589 5240
rect 893 5161 947 5413
<< metal1 >>
rect 226 5401 529 5947
rect 605 5259 686 5502
rect 605 5246 901 5259
rect 605 5175 902 5246
rect 193 3468 529 5087
rect 605 4250 686 5175
rect 978 4239 1024 5585
rect -74 3354 1232 3419
rect -74 3213 1232 3278
rect -74 3071 1232 3136
rect -74 2930 1232 2995
<< metal2 >>
rect 294 5498 529 5947
rect 294 2201 385 5249
rect 800 2189 890 3574
rect 1143 2411 1233 3757
rect 800 2096 1233 2189
<< metal3 >>
rect 4 3608 1233 3702
rect 10 3351 1270 3444
use alatch_512x8m81  alatch_512x8m81_0
timestamp 1763765945
transform 1 0 49 0 1 838
box -63 409 1197 2033
use M1_NWELL11_512x8m81  M1_NWELL11_512x8m81_0
timestamp 1763765945
transform 1 0 233 0 1 3869
box -154 -491 154 1302
use M1_POLY2$$46559276_512x8m81  M1_POLY2$$46559276_512x8m81_0
timestamp 1763765945
transform 1 0 805 0 1 5217
box -123 -48 123 48
use M1_POLY2$$46559276_512x8m81  M1_POLY2$$46559276_512x8m81_1
timestamp 1763765945
transform 1 0 448 0 1 5203
box -123 -48 123 48
use M1_PSUB$$47335468_512x8m81  M1_PSUB$$47335468_512x8m81_0
timestamp 1763765945
transform 1 0 276 0 1 5583
box -55 -190 56 400
use M2_M1$$34864172_512x8m81  M2_M1$$34864172_512x8m81_0
timestamp 1763765945
transform 1 0 413 0 1 5203
box -119 -46 119 46
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1763765945
transform 1 0 339 0 1 2322
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_1
timestamp 1763765945
transform 1 0 645 0 1 3613
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_2
timestamp 1763765945
transform 1 0 1005 0 1 4048
box -43 -122 43 122
use M2_M1$$43376684_512x8m81  M2_M1$$43376684_512x8m81_0
timestamp 1763765945
transform 1 0 853 0 1 4467
box -44 21 44 579
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_0
timestamp 1763765945
transform 1 0 339 0 1 5673
box -44 -275 44 275
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_1
timestamp 1763765945
transform 1 0 484 0 1 5673
box -44 -275 44 275
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_2
timestamp 1763765945
transform 1 0 848 0 1 5677
box -44 -275 44 275
use M2_M1$$47500332_512x8m81  M2_M1$$47500332_512x8m81_0
timestamp 1763765945
transform 1 0 493 0 1 4308
box -44 -432 44 732
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_0
timestamp 1763765945
transform 1 0 1188 0 1 3635
box -44 -123 44 123
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_1
timestamp 1763765945
transform 1 0 845 0 1 3351
box -44 -123 44 123
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_0
timestamp 1763765945
transform 1 0 339 0 1 5673
box -84 -185 84 275
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_1
timestamp 1763765945
transform 1 0 484 0 1 5673
box -84 -185 84 275
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_2
timestamp 1763765945
transform 1 0 848 0 1 5677
box -84 -185 84 275
use M3_M2$$47644716_512x8m81  M3_M2$$47644716_512x8m81_0
timestamp 1763765945
transform 1 0 493 0 1 4308
box -45 -432 45 732
use M3_M2$$47645740_512x8m81  M3_M2$$47645740_512x8m81_0
timestamp 1763765945
transform 1 0 853 0 1 4467
box -45 -579 45 579
use nmos_1p2$$47502380_512x8m81  nmos_1p2$$47502380_512x8m81_0
timestamp 1763765945
transform 1 0 907 0 1 5441
box -102 -44 130 531
use nmos_5p04310591302066_512x8m81  nmos_5p04310591302066_512x8m81_0
timestamp 1763765945
transform 1 0 525 0 1 5296
box -88 -44 144 701
use pmos_1p2$$47503404_512x8m81  pmos_1p2$$47503404_512x8m81_0
timestamp 1763765945
transform 1 0 547 0 1 3464
box -188 -86 216 1737
use pmos_1p2$$47504428_512x8m81  pmos_1p2$$47504428_512x8m81_0
timestamp 1763765945
transform 1 0 907 0 1 3899
box -188 -86 216 1314
<< end >>
