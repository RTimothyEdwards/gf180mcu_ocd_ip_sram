VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_ocd_ip_sram__sram1024x8m8wm1
  CLASS BLOCK ;
  FOREIGN gf180mcu_ocd_ip_sram__sram1024x8m8wm1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 301.300 BY 515.810 ;
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 101.520 0.000 102.305 6.000 ;
    END
  END A[8]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 103.965 0.000 104.750 6.000 ;
    END
  END A[7]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 188.200 0.000 188.985 6.000 ;
    END
  END A[6]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 190.455 0.000 191.240 6.000 ;
    END
  END A[5]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 193.070 0.000 193.855 6.000 ;
    END
  END A[4]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 196.925 0.000 197.710 6.000 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 108.005 0.000 108.790 6.000 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 113.930 0.000 114.715 6.000 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 119.850 0.000 120.630 6.000 ;
    END
  END A[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.418650 ;
    PORT
      LAYER Metal2 ;
        RECT 176.195 0.000 176.980 6.000 ;
    END
  END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.738400 ;
    PORT
      LAYER Metal2 ;
        RECT 97.775 0.000 98.560 6.000 ;
    END
  END CLK
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal1 ;
        RECT 291.455 5.200 291.795 5.265 ;
        RECT 291.230 4.800 292.020 5.200 ;
        RECT 291.455 4.735 291.795 4.800 ;
      LAYER Metal2 ;
        RECT 291.200 5.030 291.985 6.000 ;
        RECT 290.800 4.305 291.985 5.030 ;
        RECT 290.800 0.000 291.585 4.305 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal1 ;
        RECT 254.655 5.200 254.995 5.265 ;
        RECT 254.430 4.800 255.220 5.200 ;
        RECT 254.655 4.735 254.995 4.800 ;
      LAYER Metal2 ;
        RECT 254.645 5.215 254.930 6.000 ;
        RECT 254.645 4.790 254.995 5.215 ;
        RECT 254.645 4.245 254.930 4.790 ;
        RECT 254.605 0.000 255.385 4.245 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal1 ;
        RECT 249.530 5.200 249.870 5.265 ;
        RECT 249.305 4.800 250.095 5.200 ;
        RECT 249.530 4.735 249.870 4.800 ;
      LAYER Metal2 ;
        RECT 249.530 5.215 249.810 6.000 ;
        RECT 249.530 4.790 249.870 5.215 ;
        RECT 249.530 4.245 249.810 4.790 ;
        RECT 249.235 0.000 250.020 4.245 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal1 ;
        RECT 212.245 5.215 212.585 5.280 ;
        RECT 212.020 4.815 212.810 5.215 ;
        RECT 212.245 4.750 212.585 4.815 ;
      LAYER Metal2 ;
        RECT 212.255 5.230 212.625 6.000 ;
        RECT 212.245 4.805 212.625 5.230 ;
        RECT 212.255 4.355 212.625 4.805 ;
        RECT 212.255 4.350 213.940 4.355 ;
        RECT 212.255 3.985 214.845 4.350 ;
        RECT 214.060 0.000 214.845 3.985 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal1 ;
        RECT 85.695 5.260 86.035 5.325 ;
        RECT 85.470 4.860 86.260 5.260 ;
        RECT 85.695 4.795 86.035 4.860 ;
      LAYER Metal2 ;
        RECT 85.695 5.275 86.000 6.000 ;
        RECT 85.695 4.850 86.035 5.275 ;
        RECT 83.280 4.545 86.000 4.850 ;
        RECT 83.280 0.000 84.065 4.545 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal1 ;
        RECT 47.600 5.260 47.940 5.325 ;
        RECT 47.375 4.860 48.165 5.260 ;
        RECT 47.600 4.795 47.940 4.860 ;
      LAYER Metal2 ;
        RECT 48.730 5.425 49.015 6.000 ;
        RECT 47.595 5.140 49.015 5.425 ;
        RECT 47.595 4.850 47.940 5.140 ;
        RECT 47.595 4.160 47.880 4.850 ;
        RECT 47.085 3.720 47.880 4.160 ;
        RECT 47.085 0.000 47.870 3.720 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal1 ;
        RECT 43.180 5.260 43.520 5.325 ;
        RECT 42.955 4.860 43.745 5.260 ;
        RECT 43.180 4.795 43.520 4.860 ;
      LAYER Metal2 ;
        RECT 43.215 5.290 43.540 6.000 ;
        RECT 43.180 4.170 43.540 5.290 ;
        RECT 42.720 0.000 43.505 4.170 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal1 ;
        RECT 6.730 5.260 7.070 5.325 ;
        RECT 6.505 4.860 7.295 5.260 ;
        RECT 6.730 4.795 7.070 4.860 ;
      LAYER Metal2 ;
        RECT 6.520 0.000 7.305 6.000 ;
    END
  END D[0]
  PIN GWEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.141600 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal2 ;
        RECT 142.055 0.000 142.840 6.000 ;
    END
  END GWEN
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 285.870 4.245 286.200 6.000 ;
        RECT 285.490 0.000 286.275 4.245 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 257.025 4.245 257.345 6.000 ;
        RECT 256.960 0.000 257.740 4.245 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 247.175 4.245 247.460 6.000 ;
        RECT 246.880 0.000 247.665 4.245 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 217.860 4.705 218.190 6.000 ;
        RECT 217.860 4.695 220.060 4.705 ;
        RECT 217.860 4.375 220.135 4.695 ;
        RECT 219.350 0.000 220.135 4.375 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 77.980 4.130 78.315 6.000 ;
        RECT 77.975 0.000 78.760 4.130 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 51.250 5.450 51.580 6.000 ;
        RECT 49.960 5.120 51.580 5.450 ;
        RECT 49.960 4.160 50.290 5.120 ;
        RECT 49.440 3.710 50.290 4.160 ;
        RECT 49.440 0.000 50.225 3.710 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 41.545 4.725 41.875 6.000 ;
        RECT 40.840 4.395 41.875 4.725 ;
        RECT 40.840 4.200 41.170 4.395 ;
        RECT 40.365 3.555 41.170 4.200 ;
        RECT 40.365 0.000 41.145 3.555 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 12.255 5.780 12.585 6.000 ;
        RECT 12.255 5.450 14.415 5.780 ;
        RECT 14.085 4.245 14.415 5.450 ;
        RECT 13.830 0.000 14.610 4.245 ;
    END
  END Q[0]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT 103.900 509.810 194.020 510.690 ;
        RECT 7.680 5.780 25.360 6.000 ;
        RECT 29.080 5.780 64.190 6.000 ;
        RECT 29.080 5.770 46.760 5.780 ;
        RECT 67.910 5.770 85.590 6.000 ;
        RECT 212.985 5.780 230.665 6.000 ;
        RECT 234.385 5.785 269.745 6.000 ;
        RECT 234.385 5.770 252.065 5.785 ;
        RECT 273.465 5.775 291.145 6.000 ;
      LAYER Metal1 ;
        RECT 4.845 505.255 5.975 505.970 ;
        RECT 4.845 504.555 6.000 505.255 ;
        RECT 295.440 505.000 296.570 506.055 ;
        RECT 295.300 504.720 296.570 505.000 ;
        RECT 4.845 503.540 5.975 504.555 ;
        RECT 295.440 503.625 296.570 504.720 ;
        RECT 4.845 499.195 5.975 499.910 ;
        RECT 4.845 498.495 6.000 499.195 ;
        RECT 295.440 498.940 296.570 499.995 ;
        RECT 295.300 498.660 296.570 498.940 ;
        RECT 4.845 497.480 5.975 498.495 ;
        RECT 295.440 497.565 296.570 498.660 ;
        RECT 4.845 493.135 5.975 493.850 ;
        RECT 4.845 492.435 6.000 493.135 ;
        RECT 295.440 492.880 296.570 493.935 ;
        RECT 295.300 492.600 296.570 492.880 ;
        RECT 4.845 491.420 5.975 492.435 ;
        RECT 295.440 491.505 296.570 492.600 ;
        RECT 4.845 487.075 5.975 487.790 ;
        RECT 4.845 486.375 6.000 487.075 ;
        RECT 295.440 486.820 296.570 487.875 ;
        RECT 295.300 486.540 296.570 486.820 ;
        RECT 4.845 485.360 5.975 486.375 ;
        RECT 295.440 485.445 296.570 486.540 ;
        RECT 4.845 481.015 5.975 481.730 ;
        RECT 4.845 480.315 6.000 481.015 ;
        RECT 295.440 480.760 296.570 481.815 ;
        RECT 295.300 480.480 296.570 480.760 ;
        RECT 4.845 479.300 5.975 480.315 ;
        RECT 295.440 479.385 296.570 480.480 ;
        RECT 4.845 474.955 5.975 475.670 ;
        RECT 4.845 474.255 6.000 474.955 ;
        RECT 295.440 474.700 296.570 475.755 ;
        RECT 295.300 474.420 296.570 474.700 ;
        RECT 4.845 473.240 5.975 474.255 ;
        RECT 295.440 473.325 296.570 474.420 ;
        RECT 4.845 468.895 5.975 469.610 ;
        RECT 4.845 468.195 6.000 468.895 ;
        RECT 295.440 468.640 296.570 469.695 ;
        RECT 295.300 468.360 296.570 468.640 ;
        RECT 4.845 467.180 5.975 468.195 ;
        RECT 295.440 467.265 296.570 468.360 ;
        RECT 4.845 462.835 5.975 463.550 ;
        RECT 4.845 462.135 6.000 462.835 ;
        RECT 295.440 462.580 296.570 463.635 ;
        RECT 295.300 462.300 296.570 462.580 ;
        RECT 4.845 461.120 5.975 462.135 ;
        RECT 295.440 461.205 296.570 462.300 ;
        RECT 4.845 456.775 5.975 457.490 ;
        RECT 4.845 456.075 6.000 456.775 ;
        RECT 295.440 456.520 296.570 457.575 ;
        RECT 295.300 456.240 296.570 456.520 ;
        RECT 4.845 455.060 5.975 456.075 ;
        RECT 295.440 455.145 296.570 456.240 ;
        RECT 4.845 450.715 5.975 451.430 ;
        RECT 4.845 450.015 6.000 450.715 ;
        RECT 295.440 450.460 296.570 451.515 ;
        RECT 295.300 450.180 296.570 450.460 ;
        RECT 4.845 449.000 5.975 450.015 ;
        RECT 295.440 449.085 296.570 450.180 ;
        RECT 4.845 444.655 5.975 445.370 ;
        RECT 4.845 443.955 6.000 444.655 ;
        RECT 295.440 444.400 296.570 445.455 ;
        RECT 295.300 444.120 296.570 444.400 ;
        RECT 4.845 442.940 5.975 443.955 ;
        RECT 295.440 443.025 296.570 444.120 ;
        RECT 4.845 438.595 5.975 439.310 ;
        RECT 4.845 437.895 6.000 438.595 ;
        RECT 295.440 438.340 296.570 439.395 ;
        RECT 295.300 438.060 296.570 438.340 ;
        RECT 4.845 436.880 5.975 437.895 ;
        RECT 295.440 436.965 296.570 438.060 ;
        RECT 4.845 432.535 5.975 433.250 ;
        RECT 4.845 431.835 6.000 432.535 ;
        RECT 295.440 432.280 296.570 433.335 ;
        RECT 295.300 432.000 296.570 432.280 ;
        RECT 4.845 430.820 5.975 431.835 ;
        RECT 295.440 430.905 296.570 432.000 ;
        RECT 4.845 426.475 5.975 427.190 ;
        RECT 4.845 425.775 6.000 426.475 ;
        RECT 295.440 426.220 296.570 427.275 ;
        RECT 295.300 425.940 296.570 426.220 ;
        RECT 4.845 424.760 5.975 425.775 ;
        RECT 295.440 424.845 296.570 425.940 ;
        RECT 4.845 420.415 5.975 421.130 ;
        RECT 4.845 419.715 6.000 420.415 ;
        RECT 295.440 420.160 296.570 421.215 ;
        RECT 295.300 419.880 296.570 420.160 ;
        RECT 4.845 418.700 5.975 419.715 ;
        RECT 295.440 418.785 296.570 419.880 ;
        RECT 4.845 414.355 5.975 415.070 ;
        RECT 4.845 413.655 6.000 414.355 ;
        RECT 295.440 414.100 296.570 415.155 ;
        RECT 295.300 413.820 296.570 414.100 ;
        RECT 4.845 412.640 5.975 413.655 ;
        RECT 295.440 412.725 296.570 413.820 ;
        RECT 4.845 408.295 5.975 409.010 ;
        RECT 4.845 407.595 6.000 408.295 ;
        RECT 295.440 408.040 296.570 409.095 ;
        RECT 295.300 407.760 296.570 408.040 ;
        RECT 4.845 406.580 5.975 407.595 ;
        RECT 295.440 406.665 296.570 407.760 ;
        RECT 4.845 402.235 5.975 402.950 ;
        RECT 4.845 401.535 6.000 402.235 ;
        RECT 295.440 401.980 296.570 403.035 ;
        RECT 295.300 401.700 296.570 401.980 ;
        RECT 4.845 400.520 5.975 401.535 ;
        RECT 295.440 400.605 296.570 401.700 ;
        RECT 4.845 396.175 5.975 396.890 ;
        RECT 4.845 395.475 6.000 396.175 ;
        RECT 295.440 395.920 296.570 396.975 ;
        RECT 295.300 395.640 296.570 395.920 ;
        RECT 4.845 394.460 5.975 395.475 ;
        RECT 295.440 394.545 296.570 395.640 ;
        RECT 4.845 390.115 5.975 390.830 ;
        RECT 4.845 389.415 6.000 390.115 ;
        RECT 295.440 389.860 296.570 390.915 ;
        RECT 295.300 389.580 296.570 389.860 ;
        RECT 4.845 388.400 5.975 389.415 ;
        RECT 295.440 388.485 296.570 389.580 ;
        RECT 4.845 384.055 5.975 384.770 ;
        RECT 4.845 383.355 6.000 384.055 ;
        RECT 295.440 383.800 296.570 384.855 ;
        RECT 295.300 383.520 296.570 383.800 ;
        RECT 4.845 382.340 5.975 383.355 ;
        RECT 295.440 382.425 296.570 383.520 ;
        RECT 4.845 377.995 5.975 378.710 ;
        RECT 4.845 377.295 6.000 377.995 ;
        RECT 295.440 377.740 296.570 378.795 ;
        RECT 295.300 377.460 296.570 377.740 ;
        RECT 4.845 376.280 5.975 377.295 ;
        RECT 295.440 376.365 296.570 377.460 ;
        RECT 4.845 371.935 5.975 372.650 ;
        RECT 4.845 371.235 6.000 371.935 ;
        RECT 295.440 371.680 296.570 372.735 ;
        RECT 295.300 371.400 296.570 371.680 ;
        RECT 4.845 370.220 5.975 371.235 ;
        RECT 295.440 370.305 296.570 371.400 ;
        RECT 4.845 365.875 5.975 366.590 ;
        RECT 4.845 365.175 6.000 365.875 ;
        RECT 295.440 365.620 296.570 366.675 ;
        RECT 295.300 365.340 296.570 365.620 ;
        RECT 4.845 364.160 5.975 365.175 ;
        RECT 295.440 364.245 296.570 365.340 ;
        RECT 4.845 359.815 5.975 360.530 ;
        RECT 4.845 359.115 6.000 359.815 ;
        RECT 295.440 359.560 296.570 360.615 ;
        RECT 295.300 359.280 296.570 359.560 ;
        RECT 4.845 358.100 5.975 359.115 ;
        RECT 295.440 358.185 296.570 359.280 ;
        RECT 4.845 353.755 5.975 354.470 ;
        RECT 4.845 353.055 6.000 353.755 ;
        RECT 295.440 353.500 296.570 354.555 ;
        RECT 295.300 353.220 296.570 353.500 ;
        RECT 4.845 352.040 5.975 353.055 ;
        RECT 295.440 352.125 296.570 353.220 ;
        RECT 4.845 347.695 5.975 348.410 ;
        RECT 4.845 346.995 6.000 347.695 ;
        RECT 295.440 347.440 296.570 348.495 ;
        RECT 295.300 347.160 296.570 347.440 ;
        RECT 4.845 345.980 5.975 346.995 ;
        RECT 295.440 346.065 296.570 347.160 ;
        RECT 4.845 341.635 5.975 342.350 ;
        RECT 4.845 340.935 6.000 341.635 ;
        RECT 295.440 341.380 296.570 342.435 ;
        RECT 295.300 341.100 296.570 341.380 ;
        RECT 4.845 339.920 5.975 340.935 ;
        RECT 295.440 340.005 296.570 341.100 ;
        RECT 4.845 335.575 5.975 336.290 ;
        RECT 4.845 334.875 6.000 335.575 ;
        RECT 295.440 335.320 296.570 336.375 ;
        RECT 295.300 335.040 296.570 335.320 ;
        RECT 4.845 333.860 5.975 334.875 ;
        RECT 295.440 333.945 296.570 335.040 ;
        RECT 4.845 329.515 5.975 330.230 ;
        RECT 4.845 328.815 6.000 329.515 ;
        RECT 295.440 329.260 296.570 330.315 ;
        RECT 295.300 328.980 296.570 329.260 ;
        RECT 4.845 327.800 5.975 328.815 ;
        RECT 295.440 327.885 296.570 328.980 ;
        RECT 4.845 323.455 5.975 324.170 ;
        RECT 4.845 322.755 6.000 323.455 ;
        RECT 295.440 323.200 296.570 324.255 ;
        RECT 295.300 322.920 296.570 323.200 ;
        RECT 4.845 321.740 5.975 322.755 ;
        RECT 295.440 321.825 296.570 322.920 ;
        RECT 4.845 317.395 5.975 318.110 ;
        RECT 4.845 316.695 6.000 317.395 ;
        RECT 295.440 317.140 296.570 318.195 ;
        RECT 295.300 316.860 296.570 317.140 ;
        RECT 4.845 315.680 5.975 316.695 ;
        RECT 295.440 315.765 296.570 316.860 ;
        RECT 4.845 311.335 5.975 312.050 ;
        RECT 4.845 310.635 6.000 311.335 ;
        RECT 295.440 311.080 296.570 312.135 ;
        RECT 295.300 310.800 296.570 311.080 ;
        RECT 4.845 309.620 5.975 310.635 ;
        RECT 295.440 309.705 296.570 310.800 ;
        RECT 4.845 305.275 5.975 305.990 ;
        RECT 4.845 304.575 6.000 305.275 ;
        RECT 295.440 305.020 296.570 306.075 ;
        RECT 295.300 304.740 296.570 305.020 ;
        RECT 4.845 303.560 5.975 304.575 ;
        RECT 295.440 303.645 296.570 304.740 ;
        RECT 4.845 299.215 5.975 299.930 ;
        RECT 4.845 298.515 6.000 299.215 ;
        RECT 295.440 298.960 296.570 300.015 ;
        RECT 295.300 298.680 296.570 298.960 ;
        RECT 4.845 297.500 5.975 298.515 ;
        RECT 295.440 297.585 296.570 298.680 ;
        RECT 4.845 293.155 5.975 293.870 ;
        RECT 4.845 292.455 6.000 293.155 ;
        RECT 295.440 292.900 296.570 293.955 ;
        RECT 295.300 292.620 296.570 292.900 ;
        RECT 4.845 291.440 5.975 292.455 ;
        RECT 295.440 291.525 296.570 292.620 ;
        RECT 4.845 287.095 5.975 287.810 ;
        RECT 4.845 286.395 6.000 287.095 ;
        RECT 295.440 286.840 296.570 287.895 ;
        RECT 295.300 286.560 296.570 286.840 ;
        RECT 4.845 285.380 5.975 286.395 ;
        RECT 295.440 285.465 296.570 286.560 ;
        RECT 4.845 281.035 5.975 281.750 ;
        RECT 4.845 280.335 6.000 281.035 ;
        RECT 295.440 280.780 296.570 281.835 ;
        RECT 295.300 280.500 296.570 280.780 ;
        RECT 4.845 279.320 5.975 280.335 ;
        RECT 295.440 279.405 296.570 280.500 ;
        RECT 4.845 274.975 5.975 275.690 ;
        RECT 4.845 274.275 6.000 274.975 ;
        RECT 295.440 274.720 296.570 275.775 ;
        RECT 295.300 274.440 296.570 274.720 ;
        RECT 4.845 273.260 5.975 274.275 ;
        RECT 295.440 273.345 296.570 274.440 ;
        RECT 4.845 268.915 5.975 269.630 ;
        RECT 4.845 268.215 6.000 268.915 ;
        RECT 295.440 268.660 296.570 269.715 ;
        RECT 295.300 268.380 296.570 268.660 ;
        RECT 4.845 267.200 5.975 268.215 ;
        RECT 295.440 267.285 296.570 268.380 ;
        RECT 4.845 262.855 5.975 263.570 ;
        RECT 4.845 262.155 6.000 262.855 ;
        RECT 295.440 262.600 296.570 263.655 ;
        RECT 295.300 262.320 296.570 262.600 ;
        RECT 4.845 261.140 5.975 262.155 ;
        RECT 295.440 261.225 296.570 262.320 ;
        RECT 4.845 256.795 5.975 257.510 ;
        RECT 4.845 256.095 6.000 256.795 ;
        RECT 295.440 256.540 296.570 257.595 ;
        RECT 295.300 256.260 296.570 256.540 ;
        RECT 4.845 255.080 5.975 256.095 ;
        RECT 295.440 255.165 296.570 256.260 ;
        RECT 4.845 250.735 5.975 251.450 ;
        RECT 4.845 250.035 6.000 250.735 ;
        RECT 295.440 250.480 296.570 251.535 ;
        RECT 295.300 250.200 296.570 250.480 ;
        RECT 4.845 249.020 5.975 250.035 ;
        RECT 295.440 249.105 296.570 250.200 ;
        RECT 4.845 244.675 5.975 245.390 ;
        RECT 4.845 243.975 6.000 244.675 ;
        RECT 295.440 244.420 296.570 245.475 ;
        RECT 295.300 244.140 296.570 244.420 ;
        RECT 4.845 242.960 5.975 243.975 ;
        RECT 295.440 243.045 296.570 244.140 ;
        RECT 4.845 238.615 5.975 239.330 ;
        RECT 4.845 237.915 6.000 238.615 ;
        RECT 295.440 238.360 296.570 239.415 ;
        RECT 295.300 238.080 296.570 238.360 ;
        RECT 4.845 236.900 5.975 237.915 ;
        RECT 295.440 236.985 296.570 238.080 ;
        RECT 4.845 232.555 5.975 233.270 ;
        RECT 4.845 231.855 6.000 232.555 ;
        RECT 295.440 232.300 296.570 233.355 ;
        RECT 295.300 232.020 296.570 232.300 ;
        RECT 4.845 230.840 5.975 231.855 ;
        RECT 295.440 230.925 296.570 232.020 ;
        RECT 4.845 226.495 5.975 227.210 ;
        RECT 4.845 225.795 6.000 226.495 ;
        RECT 295.440 226.240 296.570 227.295 ;
        RECT 295.300 225.960 296.570 226.240 ;
        RECT 4.845 224.780 5.975 225.795 ;
        RECT 295.440 224.865 296.570 225.960 ;
        RECT 4.845 220.435 5.975 221.150 ;
        RECT 4.845 219.735 6.000 220.435 ;
        RECT 295.440 220.180 296.570 221.235 ;
        RECT 295.300 219.900 296.570 220.180 ;
        RECT 4.845 218.720 5.975 219.735 ;
        RECT 295.440 218.805 296.570 219.900 ;
        RECT 4.845 214.375 5.975 215.090 ;
        RECT 4.845 213.675 6.000 214.375 ;
        RECT 295.440 214.120 296.570 215.175 ;
        RECT 295.300 213.840 296.570 214.120 ;
        RECT 4.845 212.660 5.975 213.675 ;
        RECT 295.440 212.745 296.570 213.840 ;
        RECT 4.845 208.315 5.975 209.030 ;
        RECT 4.845 207.615 6.000 208.315 ;
        RECT 295.440 208.060 296.570 209.115 ;
        RECT 295.300 207.780 296.570 208.060 ;
        RECT 4.845 206.600 5.975 207.615 ;
        RECT 295.440 206.685 296.570 207.780 ;
        RECT 4.845 202.255 5.975 202.970 ;
        RECT 4.845 201.555 6.000 202.255 ;
        RECT 295.440 202.000 296.570 203.055 ;
        RECT 295.300 201.720 296.570 202.000 ;
        RECT 4.845 200.540 5.975 201.555 ;
        RECT 295.440 200.625 296.570 201.720 ;
        RECT 4.845 196.195 5.975 196.910 ;
        RECT 4.845 195.495 6.000 196.195 ;
        RECT 295.440 195.940 296.570 196.995 ;
        RECT 295.300 195.660 296.570 195.940 ;
        RECT 4.845 194.480 5.975 195.495 ;
        RECT 295.440 194.565 296.570 195.660 ;
        RECT 4.845 190.135 5.975 190.850 ;
        RECT 4.845 189.435 6.000 190.135 ;
        RECT 295.440 189.880 296.570 190.935 ;
        RECT 295.300 189.600 296.570 189.880 ;
        RECT 4.845 188.420 5.975 189.435 ;
        RECT 295.440 188.505 296.570 189.600 ;
        RECT 4.845 184.075 5.975 184.790 ;
        RECT 4.845 183.375 6.000 184.075 ;
        RECT 295.440 183.820 296.570 184.875 ;
        RECT 295.300 183.540 296.570 183.820 ;
        RECT 4.845 182.360 5.975 183.375 ;
        RECT 295.440 182.445 296.570 183.540 ;
        RECT 4.845 178.015 5.975 178.730 ;
        RECT 4.845 177.315 6.000 178.015 ;
        RECT 295.440 177.760 296.570 178.815 ;
        RECT 295.300 177.480 296.570 177.760 ;
        RECT 4.845 176.300 5.975 177.315 ;
        RECT 295.440 176.385 296.570 177.480 ;
        RECT 4.845 171.955 5.975 172.670 ;
        RECT 4.845 171.255 6.000 171.955 ;
        RECT 295.440 171.700 296.570 172.755 ;
        RECT 295.300 171.420 296.570 171.700 ;
        RECT 4.845 170.240 5.975 171.255 ;
        RECT 295.440 170.325 296.570 171.420 ;
        RECT 4.845 165.895 5.975 166.610 ;
        RECT 4.845 165.195 6.000 165.895 ;
        RECT 295.440 165.640 296.570 166.695 ;
        RECT 295.300 165.360 296.570 165.640 ;
        RECT 4.845 164.180 5.975 165.195 ;
        RECT 295.440 164.265 296.570 165.360 ;
        RECT 4.845 159.835 5.975 160.550 ;
        RECT 4.845 159.135 6.000 159.835 ;
        RECT 295.440 159.580 296.570 160.635 ;
        RECT 295.300 159.300 296.570 159.580 ;
        RECT 4.845 158.120 5.975 159.135 ;
        RECT 295.440 158.205 296.570 159.300 ;
        RECT 4.845 153.775 5.975 154.490 ;
        RECT 4.845 153.075 6.000 153.775 ;
        RECT 295.440 153.520 296.570 154.575 ;
        RECT 295.300 153.240 296.570 153.520 ;
        RECT 4.845 152.060 5.975 153.075 ;
        RECT 295.440 152.145 296.570 153.240 ;
        RECT 4.845 147.715 5.975 148.430 ;
        RECT 4.845 147.015 6.000 147.715 ;
        RECT 295.440 147.460 296.570 148.515 ;
        RECT 295.300 147.180 296.570 147.460 ;
        RECT 4.845 146.000 5.975 147.015 ;
        RECT 295.440 146.085 296.570 147.180 ;
        RECT 4.845 141.655 5.975 142.370 ;
        RECT 4.845 140.955 6.000 141.655 ;
        RECT 295.440 141.400 296.570 142.455 ;
        RECT 295.300 141.120 296.570 141.400 ;
        RECT 4.845 139.940 5.975 140.955 ;
        RECT 295.440 140.025 296.570 141.120 ;
        RECT 4.845 135.595 5.975 136.310 ;
        RECT 4.845 134.895 6.000 135.595 ;
        RECT 295.440 135.340 296.570 136.395 ;
        RECT 295.300 135.060 296.570 135.340 ;
        RECT 4.845 133.880 5.975 134.895 ;
        RECT 295.440 133.965 296.570 135.060 ;
        RECT 4.845 129.535 5.975 130.250 ;
        RECT 4.845 128.835 6.000 129.535 ;
        RECT 295.440 129.280 296.570 130.335 ;
        RECT 295.300 129.000 296.570 129.280 ;
        RECT 4.845 127.820 5.975 128.835 ;
        RECT 295.440 127.905 296.570 129.000 ;
        RECT 4.845 123.475 5.975 124.190 ;
        RECT 4.845 122.775 6.000 123.475 ;
        RECT 295.440 123.220 296.570 124.275 ;
        RECT 295.300 122.940 296.570 123.220 ;
        RECT 4.845 121.760 5.975 122.775 ;
        RECT 295.440 121.845 296.570 122.940 ;
        RECT 4.845 117.415 5.975 118.130 ;
        RECT 4.845 116.715 6.000 117.415 ;
        RECT 295.440 117.160 296.570 118.215 ;
        RECT 295.300 116.880 296.570 117.160 ;
        RECT 4.845 115.700 5.975 116.715 ;
        RECT 295.440 115.785 296.570 116.880 ;
        RECT 93.700 5.990 95.245 6.000 ;
      LAYER Metal2 ;
        RECT 2.470 512.860 298.830 513.010 ;
        RECT 2.465 509.810 298.830 512.860 ;
        RECT 2.465 509.510 6.000 509.810 ;
        RECT 295.300 509.510 298.830 509.810 ;
        RECT 2.465 505.970 5.970 509.510 ;
        RECT 295.445 506.055 298.830 509.510 ;
        RECT 2.465 503.540 5.975 505.970 ;
        RECT 295.440 503.625 298.830 506.055 ;
        RECT 2.465 499.910 5.970 503.540 ;
        RECT 295.445 499.995 298.830 503.625 ;
        RECT 2.465 497.480 5.975 499.910 ;
        RECT 295.440 497.565 298.830 499.995 ;
        RECT 2.465 493.850 5.970 497.480 ;
        RECT 295.445 493.935 298.830 497.565 ;
        RECT 2.465 491.420 5.975 493.850 ;
        RECT 295.440 491.505 298.830 493.935 ;
        RECT 2.465 487.790 5.970 491.420 ;
        RECT 295.445 487.875 298.830 491.505 ;
        RECT 2.465 485.360 5.975 487.790 ;
        RECT 295.440 485.445 298.830 487.875 ;
        RECT 2.465 481.730 5.970 485.360 ;
        RECT 295.445 481.815 298.830 485.445 ;
        RECT 2.465 479.300 5.975 481.730 ;
        RECT 295.440 479.385 298.830 481.815 ;
        RECT 2.465 475.670 5.970 479.300 ;
        RECT 295.445 475.755 298.830 479.385 ;
        RECT 2.465 473.240 5.975 475.670 ;
        RECT 295.440 473.325 298.830 475.755 ;
        RECT 2.465 469.610 5.970 473.240 ;
        RECT 295.445 469.695 298.830 473.325 ;
        RECT 2.465 467.180 5.975 469.610 ;
        RECT 295.440 467.265 298.830 469.695 ;
        RECT 2.465 463.550 5.970 467.180 ;
        RECT 295.445 463.635 298.830 467.265 ;
        RECT 2.465 461.120 5.975 463.550 ;
        RECT 295.440 461.205 298.830 463.635 ;
        RECT 2.465 457.490 5.970 461.120 ;
        RECT 295.445 457.575 298.830 461.205 ;
        RECT 2.465 455.060 5.975 457.490 ;
        RECT 295.440 455.145 298.830 457.575 ;
        RECT 2.465 451.430 5.970 455.060 ;
        RECT 295.445 451.515 298.830 455.145 ;
        RECT 2.465 449.000 5.975 451.430 ;
        RECT 295.440 449.085 298.830 451.515 ;
        RECT 2.465 445.370 5.970 449.000 ;
        RECT 295.445 445.455 298.830 449.085 ;
        RECT 2.465 442.940 5.975 445.370 ;
        RECT 295.440 443.025 298.830 445.455 ;
        RECT 2.465 439.310 5.970 442.940 ;
        RECT 295.445 439.395 298.830 443.025 ;
        RECT 2.465 436.880 5.975 439.310 ;
        RECT 295.440 436.965 298.830 439.395 ;
        RECT 2.465 433.250 5.970 436.880 ;
        RECT 295.445 433.335 298.830 436.965 ;
        RECT 2.465 430.820 5.975 433.250 ;
        RECT 295.440 430.905 298.830 433.335 ;
        RECT 2.465 427.190 5.970 430.820 ;
        RECT 295.445 427.275 298.830 430.905 ;
        RECT 2.465 424.760 5.975 427.190 ;
        RECT 295.440 424.845 298.830 427.275 ;
        RECT 2.465 421.130 5.970 424.760 ;
        RECT 295.445 421.215 298.830 424.845 ;
        RECT 2.465 418.700 5.975 421.130 ;
        RECT 295.440 418.785 298.830 421.215 ;
        RECT 2.465 415.070 5.970 418.700 ;
        RECT 295.445 415.155 298.830 418.785 ;
        RECT 2.465 412.640 5.975 415.070 ;
        RECT 295.440 412.725 298.830 415.155 ;
        RECT 2.465 409.010 5.970 412.640 ;
        RECT 295.445 409.095 298.830 412.725 ;
        RECT 2.465 406.580 5.975 409.010 ;
        RECT 295.440 406.665 298.830 409.095 ;
        RECT 2.465 402.950 5.970 406.580 ;
        RECT 295.445 403.035 298.830 406.665 ;
        RECT 2.465 400.520 5.975 402.950 ;
        RECT 295.440 400.605 298.830 403.035 ;
        RECT 2.465 396.890 5.970 400.520 ;
        RECT 295.445 396.975 298.830 400.605 ;
        RECT 2.465 394.460 5.975 396.890 ;
        RECT 295.440 394.545 298.830 396.975 ;
        RECT 2.465 390.830 5.970 394.460 ;
        RECT 295.445 390.915 298.830 394.545 ;
        RECT 2.465 388.400 5.975 390.830 ;
        RECT 295.440 388.485 298.830 390.915 ;
        RECT 2.465 384.770 5.970 388.400 ;
        RECT 295.445 384.855 298.830 388.485 ;
        RECT 2.465 382.340 5.975 384.770 ;
        RECT 295.440 382.425 298.830 384.855 ;
        RECT 2.465 378.710 5.970 382.340 ;
        RECT 295.445 378.795 298.830 382.425 ;
        RECT 2.465 376.280 5.975 378.710 ;
        RECT 295.440 376.365 298.830 378.795 ;
        RECT 2.465 372.650 5.970 376.280 ;
        RECT 295.445 372.735 298.830 376.365 ;
        RECT 2.465 370.220 5.975 372.650 ;
        RECT 295.440 370.305 298.830 372.735 ;
        RECT 2.465 366.590 5.970 370.220 ;
        RECT 295.445 366.675 298.830 370.305 ;
        RECT 2.465 364.160 5.975 366.590 ;
        RECT 295.440 364.245 298.830 366.675 ;
        RECT 2.465 360.530 5.970 364.160 ;
        RECT 295.445 360.615 298.830 364.245 ;
        RECT 2.465 358.100 5.975 360.530 ;
        RECT 295.440 358.185 298.830 360.615 ;
        RECT 2.465 354.470 5.970 358.100 ;
        RECT 295.445 354.555 298.830 358.185 ;
        RECT 2.465 352.040 5.975 354.470 ;
        RECT 295.440 352.125 298.830 354.555 ;
        RECT 2.465 348.410 5.970 352.040 ;
        RECT 295.445 348.495 298.830 352.125 ;
        RECT 2.465 345.980 5.975 348.410 ;
        RECT 295.440 346.065 298.830 348.495 ;
        RECT 2.465 342.350 5.970 345.980 ;
        RECT 295.445 342.435 298.830 346.065 ;
        RECT 2.465 339.920 5.975 342.350 ;
        RECT 295.440 340.005 298.830 342.435 ;
        RECT 2.465 336.290 5.970 339.920 ;
        RECT 295.445 336.375 298.830 340.005 ;
        RECT 2.465 333.860 5.975 336.290 ;
        RECT 295.440 333.945 298.830 336.375 ;
        RECT 2.465 330.230 5.970 333.860 ;
        RECT 295.445 330.315 298.830 333.945 ;
        RECT 2.465 327.800 5.975 330.230 ;
        RECT 295.440 327.885 298.830 330.315 ;
        RECT 2.465 324.170 5.970 327.800 ;
        RECT 295.445 324.255 298.830 327.885 ;
        RECT 2.465 321.740 5.975 324.170 ;
        RECT 295.440 321.825 298.830 324.255 ;
        RECT 2.465 318.110 5.970 321.740 ;
        RECT 295.445 318.195 298.830 321.825 ;
        RECT 2.465 315.680 5.975 318.110 ;
        RECT 295.440 315.765 298.830 318.195 ;
        RECT 2.465 312.050 5.970 315.680 ;
        RECT 295.445 312.270 298.830 315.765 ;
        RECT 2.465 309.620 5.975 312.050 ;
        RECT 2.465 305.990 5.970 309.620 ;
        RECT 2.465 303.560 5.975 305.990 ;
        RECT 2.465 299.930 5.970 303.560 ;
        RECT 2.465 297.500 5.975 299.930 ;
        RECT 2.465 293.870 5.970 297.500 ;
        RECT 2.465 291.440 5.975 293.870 ;
        RECT 2.465 287.810 5.970 291.440 ;
        RECT 2.465 285.380 5.975 287.810 ;
        RECT 2.465 281.750 5.970 285.380 ;
        RECT 2.465 279.320 5.975 281.750 ;
        RECT 2.465 275.690 5.970 279.320 ;
        RECT 2.465 273.260 5.975 275.690 ;
        RECT 2.465 269.630 5.970 273.260 ;
        RECT 2.465 267.200 5.975 269.630 ;
        RECT 2.465 263.570 5.970 267.200 ;
        RECT 2.465 261.140 5.975 263.570 ;
        RECT 2.465 257.510 5.970 261.140 ;
        RECT 2.465 255.080 5.975 257.510 ;
        RECT 2.465 251.450 5.970 255.080 ;
        RECT 2.465 249.020 5.975 251.450 ;
        RECT 2.465 245.390 5.970 249.020 ;
        RECT 2.465 242.960 5.975 245.390 ;
        RECT 2.465 239.330 5.970 242.960 ;
        RECT 2.465 236.900 5.975 239.330 ;
        RECT 2.465 233.270 5.970 236.900 ;
        RECT 2.465 230.840 5.975 233.270 ;
        RECT 2.465 227.210 5.970 230.840 ;
        RECT 2.465 224.780 5.975 227.210 ;
        RECT 2.465 221.150 5.970 224.780 ;
        RECT 2.465 218.720 5.975 221.150 ;
        RECT 2.465 215.090 5.970 218.720 ;
        RECT 2.465 212.660 5.975 215.090 ;
        RECT 2.465 209.030 5.970 212.660 ;
        RECT 2.465 206.600 5.975 209.030 ;
        RECT 2.465 202.970 5.970 206.600 ;
        RECT 2.465 200.540 5.975 202.970 ;
        RECT 2.465 196.910 5.970 200.540 ;
        RECT 2.465 194.480 5.975 196.910 ;
        RECT 2.465 190.850 5.970 194.480 ;
        RECT 2.465 188.420 5.975 190.850 ;
        RECT 2.465 184.790 5.970 188.420 ;
        RECT 2.465 182.360 5.975 184.790 ;
        RECT 2.465 178.730 5.970 182.360 ;
        RECT 2.465 176.300 5.975 178.730 ;
        RECT 2.465 172.670 5.970 176.300 ;
        RECT 2.465 170.240 5.975 172.670 ;
        RECT 2.465 166.610 5.970 170.240 ;
        RECT 295.440 168.360 298.830 312.270 ;
        RECT 2.465 164.180 5.975 166.610 ;
        RECT 2.465 160.550 5.970 164.180 ;
        RECT 2.465 158.120 5.975 160.550 ;
        RECT 2.465 154.490 5.970 158.120 ;
        RECT 2.465 152.060 5.975 154.490 ;
        RECT 2.465 148.430 5.970 152.060 ;
        RECT 2.465 146.000 5.975 148.430 ;
        RECT 2.465 142.370 5.970 146.000 ;
        RECT 2.465 139.940 5.975 142.370 ;
        RECT 2.465 136.310 5.970 139.940 ;
        RECT 2.465 133.880 5.975 136.310 ;
        RECT 2.465 130.250 5.970 133.880 ;
        RECT 2.465 127.820 5.975 130.250 ;
        RECT 2.465 124.190 5.970 127.820 ;
        RECT 2.465 121.760 5.975 124.190 ;
        RECT 2.465 118.130 5.970 121.760 ;
        RECT 2.465 115.700 5.975 118.130 ;
        RECT 2.465 110.435 5.970 115.700 ;
        RECT 295.440 110.435 298.835 168.360 ;
        RECT 2.465 4.330 5.975 110.435 ;
        RECT 26.795 4.830 27.580 6.000 ;
        RECT 65.605 4.830 66.390 6.000 ;
        RECT 2.465 1.410 5.970 4.330 ;
        RECT 88.750 4.285 89.535 6.000 ;
        RECT 93.695 5.965 95.245 6.000 ;
        RECT 131.250 5.180 132.035 6.000 ;
        RECT 137.620 5.180 138.405 6.000 ;
        RECT 207.850 4.315 208.635 6.000 ;
        RECT 232.070 4.830 232.855 6.000 ;
        RECT 271.220 4.810 272.005 6.000 ;
        RECT 295.330 4.330 298.835 110.435 ;
        RECT 2.470 0.985 5.970 1.410 ;
        RECT 295.330 0.985 298.830 4.330 ;
      LAYER Metal3 ;
        RECT 5.090 513.680 8.590 515.810 ;
        RECT 5.090 513.010 8.585 513.680 ;
        RECT 14.480 513.010 17.975 515.810 ;
        RECT 24.630 513.680 28.130 515.810 ;
        RECT 33.380 515.110 36.880 515.810 ;
        RECT 24.630 513.010 28.125 513.680 ;
        RECT 33.380 513.010 36.875 515.110 ;
        RECT 44.170 513.010 47.665 515.810 ;
        RECT 52.280 513.010 55.775 515.810 ;
        RECT 63.710 513.010 67.205 515.810 ;
        RECT 72.285 513.010 75.780 515.810 ;
        RECT 84.680 513.680 88.180 515.810 ;
        RECT 84.685 513.010 88.180 513.680 ;
        RECT 93.000 513.010 96.495 515.810 ;
        RECT 107.485 513.010 110.980 515.810 ;
        RECT 123.950 513.010 127.445 515.810 ;
        RECT 135.045 513.010 138.540 515.810 ;
        RECT 144.305 513.010 147.800 515.810 ;
        RECT 157.740 513.010 161.235 515.810 ;
        RECT 162.095 513.010 165.590 515.810 ;
        RECT 171.155 513.010 174.650 515.810 ;
        RECT 183.990 513.010 187.485 515.810 ;
        RECT 189.915 513.010 193.410 515.810 ;
        RECT 201.415 513.010 204.910 515.810 ;
        RECT 210.520 513.010 214.015 515.810 ;
        RECT 221.995 513.010 225.490 515.810 ;
        RECT 230.060 513.010 233.555 515.810 ;
        RECT 240.895 513.010 244.390 515.810 ;
        RECT 249.600 513.010 253.095 515.810 ;
        RECT 259.795 513.010 263.290 515.810 ;
        RECT 269.125 513.010 272.620 515.810 ;
        RECT 279.300 513.010 282.795 515.810 ;
        RECT 290.115 513.010 293.610 515.810 ;
        RECT 295.330 513.010 298.825 515.810 ;
        RECT 0.000 509.810 301.300 513.010 ;
        RECT 0.000 509.510 6.000 509.810 ;
        RECT 295.300 509.510 301.300 509.810 ;
        RECT 5.090 509.505 6.000 509.510 ;
        RECT 296.440 506.055 301.300 506.065 ;
        RECT 0.000 503.530 5.975 505.980 ;
        RECT 295.440 503.625 301.300 506.055 ;
        RECT 296.440 503.615 301.300 503.625 ;
        RECT 296.440 499.995 301.300 500.005 ;
        RECT 0.000 497.470 5.975 499.920 ;
        RECT 295.440 497.565 301.300 499.995 ;
        RECT 296.440 497.555 301.300 497.565 ;
        RECT 296.440 493.935 301.300 493.945 ;
        RECT 0.000 491.410 5.975 493.860 ;
        RECT 295.440 491.505 301.300 493.935 ;
        RECT 296.440 491.495 301.300 491.505 ;
        RECT 296.440 487.875 301.300 487.885 ;
        RECT 0.000 485.350 5.975 487.800 ;
        RECT 295.440 485.445 301.300 487.875 ;
        RECT 296.440 485.435 301.300 485.445 ;
        RECT 296.440 481.815 301.300 481.825 ;
        RECT 0.000 479.290 5.975 481.740 ;
        RECT 295.440 479.385 301.300 481.815 ;
        RECT 296.440 479.375 301.300 479.385 ;
        RECT 296.440 475.755 301.300 475.765 ;
        RECT 0.000 473.230 5.975 475.680 ;
        RECT 295.440 473.325 301.300 475.755 ;
        RECT 296.440 473.315 301.300 473.325 ;
        RECT 296.440 469.695 301.300 469.705 ;
        RECT 0.000 467.170 5.975 469.620 ;
        RECT 295.440 467.265 301.300 469.695 ;
        RECT 296.440 467.255 301.300 467.265 ;
        RECT 296.440 463.635 301.300 463.645 ;
        RECT 0.000 461.110 5.975 463.560 ;
        RECT 295.440 461.205 301.300 463.635 ;
        RECT 296.440 461.195 301.300 461.205 ;
        RECT 296.440 457.575 301.300 457.585 ;
        RECT 0.000 455.050 5.975 457.500 ;
        RECT 295.440 455.145 301.300 457.575 ;
        RECT 296.440 455.135 301.300 455.145 ;
        RECT 296.440 451.515 301.300 451.525 ;
        RECT 0.000 448.990 5.975 451.440 ;
        RECT 295.440 449.085 301.300 451.515 ;
        RECT 296.440 449.075 301.300 449.085 ;
        RECT 296.440 445.455 301.300 445.465 ;
        RECT 0.000 442.930 5.975 445.380 ;
        RECT 295.440 443.025 301.300 445.455 ;
        RECT 296.440 443.015 301.300 443.025 ;
        RECT 296.440 439.395 301.300 439.405 ;
        RECT 0.000 436.870 5.975 439.320 ;
        RECT 295.440 436.965 301.300 439.395 ;
        RECT 296.440 436.955 301.300 436.965 ;
        RECT 296.440 433.335 301.300 433.345 ;
        RECT 0.000 430.810 5.975 433.260 ;
        RECT 295.440 430.905 301.300 433.335 ;
        RECT 296.440 430.895 301.300 430.905 ;
        RECT 296.440 427.275 301.300 427.285 ;
        RECT 0.000 424.750 5.975 427.200 ;
        RECT 295.440 424.845 301.300 427.275 ;
        RECT 296.440 424.835 301.300 424.845 ;
        RECT 296.440 421.215 301.300 421.225 ;
        RECT 0.000 418.690 5.975 421.140 ;
        RECT 295.440 418.785 301.300 421.215 ;
        RECT 296.440 418.775 301.300 418.785 ;
        RECT 296.440 415.155 301.300 415.165 ;
        RECT 0.000 412.630 5.975 415.080 ;
        RECT 295.440 412.725 301.300 415.155 ;
        RECT 296.440 412.715 301.300 412.725 ;
        RECT 296.440 409.095 301.300 409.105 ;
        RECT 0.000 406.570 5.975 409.020 ;
        RECT 295.440 406.665 301.300 409.095 ;
        RECT 296.440 406.655 301.300 406.665 ;
        RECT 296.440 403.035 301.300 403.045 ;
        RECT 0.000 400.510 5.975 402.960 ;
        RECT 295.440 400.605 301.300 403.035 ;
        RECT 296.440 400.595 301.300 400.605 ;
        RECT 296.440 396.975 301.300 396.985 ;
        RECT 0.000 394.450 5.975 396.900 ;
        RECT 295.440 394.545 301.300 396.975 ;
        RECT 296.440 394.535 301.300 394.545 ;
        RECT 296.440 390.915 301.300 390.925 ;
        RECT 0.000 388.390 5.975 390.840 ;
        RECT 295.440 388.485 301.300 390.915 ;
        RECT 296.440 388.475 301.300 388.485 ;
        RECT 296.440 384.855 301.300 384.865 ;
        RECT 0.000 382.330 5.975 384.780 ;
        RECT 295.440 382.425 301.300 384.855 ;
        RECT 296.440 382.415 301.300 382.425 ;
        RECT 296.440 378.795 301.300 378.805 ;
        RECT 0.000 376.270 5.975 378.720 ;
        RECT 295.440 376.365 301.300 378.795 ;
        RECT 296.440 376.355 301.300 376.365 ;
        RECT 296.440 372.735 301.300 372.745 ;
        RECT 0.000 370.210 5.975 372.660 ;
        RECT 295.440 370.305 301.300 372.735 ;
        RECT 296.440 370.295 301.300 370.305 ;
        RECT 296.440 366.675 301.300 366.685 ;
        RECT 0.000 364.150 5.975 366.600 ;
        RECT 295.440 364.245 301.300 366.675 ;
        RECT 296.440 364.235 301.300 364.245 ;
        RECT 296.440 360.615 301.300 360.625 ;
        RECT 0.000 358.090 5.975 360.540 ;
        RECT 295.440 358.185 301.300 360.615 ;
        RECT 296.440 358.175 301.300 358.185 ;
        RECT 296.440 354.555 301.300 354.565 ;
        RECT 0.000 352.030 5.975 354.480 ;
        RECT 295.440 352.125 301.300 354.555 ;
        RECT 296.440 352.115 301.300 352.125 ;
        RECT 296.440 348.495 301.300 348.505 ;
        RECT 0.000 345.970 5.975 348.420 ;
        RECT 295.440 346.065 301.300 348.495 ;
        RECT 296.440 346.055 301.300 346.065 ;
        RECT 296.440 342.435 301.300 342.445 ;
        RECT 0.000 339.910 5.975 342.360 ;
        RECT 295.440 340.005 301.300 342.435 ;
        RECT 296.440 339.995 301.300 340.005 ;
        RECT 296.440 336.375 301.300 336.385 ;
        RECT 0.000 333.850 5.975 336.300 ;
        RECT 295.440 333.945 301.300 336.375 ;
        RECT 296.440 333.935 301.300 333.945 ;
        RECT 296.440 330.315 301.300 330.325 ;
        RECT 0.000 327.790 5.975 330.240 ;
        RECT 295.440 327.885 301.300 330.315 ;
        RECT 296.440 327.875 301.300 327.885 ;
        RECT 296.440 324.255 301.300 324.265 ;
        RECT 0.000 321.730 5.975 324.180 ;
        RECT 295.440 321.825 301.300 324.255 ;
        RECT 296.440 321.815 301.300 321.825 ;
        RECT 296.440 318.195 301.300 318.205 ;
        RECT 0.000 315.670 5.975 318.120 ;
        RECT 295.440 315.765 301.300 318.195 ;
        RECT 296.440 315.755 301.300 315.765 ;
        RECT 296.440 312.135 301.300 312.145 ;
        RECT 0.000 309.610 5.975 312.060 ;
        RECT 295.440 309.705 301.300 312.135 ;
        RECT 296.440 309.695 301.300 309.705 ;
        RECT 296.440 306.075 301.300 306.085 ;
        RECT 0.000 303.550 5.975 306.000 ;
        RECT 295.440 303.645 301.300 306.075 ;
        RECT 296.440 303.635 301.300 303.645 ;
        RECT 296.440 300.015 301.300 300.025 ;
        RECT 0.000 297.490 5.975 299.940 ;
        RECT 295.440 297.585 301.300 300.015 ;
        RECT 296.440 297.575 301.300 297.585 ;
        RECT 296.440 293.955 301.300 293.965 ;
        RECT 0.000 291.430 5.975 293.880 ;
        RECT 295.440 291.525 301.300 293.955 ;
        RECT 296.440 291.515 301.300 291.525 ;
        RECT 296.440 287.895 301.300 287.905 ;
        RECT 0.000 285.370 5.975 287.820 ;
        RECT 295.440 285.465 301.300 287.895 ;
        RECT 296.440 285.455 301.300 285.465 ;
        RECT 296.440 281.835 301.300 281.845 ;
        RECT 0.000 279.310 5.975 281.760 ;
        RECT 295.440 279.405 301.300 281.835 ;
        RECT 296.440 279.395 301.300 279.405 ;
        RECT 296.440 275.775 301.300 275.785 ;
        RECT 0.000 273.250 5.975 275.700 ;
        RECT 295.440 273.345 301.300 275.775 ;
        RECT 296.440 273.335 301.300 273.345 ;
        RECT 296.440 269.715 301.300 269.725 ;
        RECT 0.000 267.190 5.975 269.640 ;
        RECT 295.440 267.285 301.300 269.715 ;
        RECT 296.440 267.275 301.300 267.285 ;
        RECT 296.440 263.655 301.300 263.665 ;
        RECT 0.000 261.130 5.975 263.580 ;
        RECT 295.440 261.225 301.300 263.655 ;
        RECT 296.440 261.215 301.300 261.225 ;
        RECT 296.440 257.595 301.300 257.605 ;
        RECT 0.000 255.070 5.975 257.520 ;
        RECT 295.440 255.165 301.300 257.595 ;
        RECT 296.440 255.155 301.300 255.165 ;
        RECT 296.440 251.535 301.300 251.545 ;
        RECT 0.000 249.010 5.975 251.460 ;
        RECT 295.440 249.105 301.300 251.535 ;
        RECT 296.440 249.095 301.300 249.105 ;
        RECT 296.440 245.475 301.300 245.485 ;
        RECT 0.000 242.950 5.975 245.400 ;
        RECT 295.440 243.045 301.300 245.475 ;
        RECT 296.440 243.035 301.300 243.045 ;
        RECT 296.440 239.415 301.300 239.425 ;
        RECT 0.000 236.890 5.975 239.340 ;
        RECT 295.440 236.985 301.300 239.415 ;
        RECT 296.440 236.975 301.300 236.985 ;
        RECT 296.440 233.355 301.300 233.365 ;
        RECT 0.000 230.830 5.975 233.280 ;
        RECT 295.440 230.925 301.300 233.355 ;
        RECT 296.440 230.915 301.300 230.925 ;
        RECT 296.440 227.295 301.300 227.305 ;
        RECT 0.000 224.770 5.975 227.220 ;
        RECT 295.440 224.865 301.300 227.295 ;
        RECT 296.440 224.855 301.300 224.865 ;
        RECT 296.440 221.235 301.300 221.245 ;
        RECT 0.000 218.710 5.975 221.160 ;
        RECT 295.440 218.805 301.300 221.235 ;
        RECT 296.440 218.795 301.300 218.805 ;
        RECT 296.440 215.175 301.300 215.185 ;
        RECT 0.000 212.650 5.975 215.100 ;
        RECT 295.440 212.745 301.300 215.175 ;
        RECT 296.440 212.735 301.300 212.745 ;
        RECT 296.440 209.115 301.300 209.125 ;
        RECT 0.000 206.590 5.975 209.040 ;
        RECT 295.440 206.685 301.300 209.115 ;
        RECT 296.440 206.675 301.300 206.685 ;
        RECT 296.440 203.055 301.300 203.065 ;
        RECT 0.000 200.530 5.975 202.980 ;
        RECT 295.440 200.625 301.300 203.055 ;
        RECT 296.440 200.615 301.300 200.625 ;
        RECT 296.440 196.995 301.300 197.005 ;
        RECT 0.000 194.470 5.975 196.920 ;
        RECT 295.440 194.565 301.300 196.995 ;
        RECT 296.440 194.555 301.300 194.565 ;
        RECT 296.440 190.935 301.300 190.945 ;
        RECT 0.000 188.410 5.975 190.860 ;
        RECT 295.440 188.505 301.300 190.935 ;
        RECT 296.440 188.495 301.300 188.505 ;
        RECT 296.440 184.875 301.300 184.885 ;
        RECT 0.000 182.350 5.975 184.800 ;
        RECT 295.440 182.445 301.300 184.875 ;
        RECT 296.440 182.435 301.300 182.445 ;
        RECT 296.440 178.815 301.300 178.825 ;
        RECT 0.000 176.290 5.975 178.740 ;
        RECT 295.440 176.385 301.300 178.815 ;
        RECT 296.440 176.375 301.300 176.385 ;
        RECT 296.440 172.755 301.300 172.765 ;
        RECT 0.000 170.230 5.975 172.680 ;
        RECT 295.440 170.325 301.300 172.755 ;
        RECT 296.440 170.315 301.300 170.325 ;
        RECT 296.440 166.695 301.300 166.705 ;
        RECT 0.000 164.170 5.975 166.620 ;
        RECT 295.440 164.265 301.300 166.695 ;
        RECT 296.440 164.255 301.300 164.265 ;
        RECT 296.440 160.635 301.300 160.645 ;
        RECT 0.000 158.110 5.975 160.560 ;
        RECT 295.440 158.205 301.300 160.635 ;
        RECT 296.440 158.195 301.300 158.205 ;
        RECT 296.440 154.575 301.300 154.585 ;
        RECT 0.000 152.050 5.975 154.500 ;
        RECT 295.440 152.145 301.300 154.575 ;
        RECT 296.440 152.135 301.300 152.145 ;
        RECT 296.440 148.515 301.300 148.525 ;
        RECT 0.000 145.990 5.975 148.440 ;
        RECT 295.440 146.085 301.300 148.515 ;
        RECT 296.440 146.075 301.300 146.085 ;
        RECT 296.440 142.455 301.300 142.465 ;
        RECT 0.000 139.930 5.975 142.380 ;
        RECT 295.440 140.025 301.300 142.455 ;
        RECT 296.440 140.015 301.300 140.025 ;
        RECT 296.440 136.395 301.300 136.405 ;
        RECT 0.000 133.870 5.975 136.320 ;
        RECT 295.440 133.965 301.300 136.395 ;
        RECT 296.440 133.955 301.300 133.965 ;
        RECT 296.440 130.335 301.300 130.345 ;
        RECT 0.000 127.810 5.975 130.260 ;
        RECT 295.440 127.905 301.300 130.335 ;
        RECT 296.440 127.895 301.300 127.905 ;
        RECT 296.440 124.275 301.300 124.285 ;
        RECT 0.000 121.750 5.975 124.200 ;
        RECT 295.440 121.845 301.300 124.275 ;
        RECT 296.440 121.835 301.300 121.845 ;
        RECT 296.440 118.215 301.300 118.225 ;
        RECT 0.000 115.690 5.975 118.140 ;
        RECT 295.440 115.785 301.300 118.215 ;
        RECT 296.440 115.775 301.300 115.785 ;
        RECT 0.000 109.905 3.545 109.910 ;
        RECT 297.750 109.905 301.300 109.910 ;
        RECT 0.000 102.880 6.000 109.905 ;
        RECT 295.300 102.880 301.300 109.905 ;
        RECT 0.000 96.170 5.975 102.880 ;
        RECT 295.335 96.170 301.300 102.880 ;
        RECT 0.000 95.175 6.000 96.170 ;
        RECT 295.300 95.175 301.300 96.170 ;
        RECT 300.600 95.170 301.300 95.175 ;
        RECT 295.300 85.600 295.500 86.350 ;
        RECT 295.300 84.370 295.500 85.125 ;
        RECT 0.000 78.350 3.545 78.355 ;
        RECT 297.750 78.350 301.300 78.355 ;
        RECT 0.000 76.400 5.975 78.350 ;
        RECT 295.335 76.400 301.300 78.350 ;
        RECT 0.000 74.855 6.000 76.400 ;
        RECT 0.010 74.850 6.000 74.855 ;
        RECT 295.300 74.850 301.300 76.400 ;
        RECT 297.750 67.740 301.300 67.750 ;
        RECT 0.010 67.735 6.000 67.740 ;
        RECT 0.000 58.210 6.000 67.735 ;
        RECT 295.300 58.210 301.300 67.740 ;
        RECT 0.000 58.205 0.700 58.210 ;
        RECT 300.600 58.205 301.300 58.210 ;
        RECT 0.000 47.315 3.545 47.325 ;
        RECT 300.600 47.315 301.300 47.320 ;
        RECT 0.000 44.810 6.000 47.315 ;
        RECT 295.300 44.810 301.300 47.315 ;
        RECT 0.000 42.955 5.975 44.810 ;
        RECT 295.335 42.970 301.300 44.810 ;
        RECT 0.000 40.125 6.000 42.955 ;
        RECT 0.010 40.120 6.000 40.125 ;
        RECT 295.300 40.120 301.300 42.970 ;
        RECT 0.010 40.020 5.975 40.120 ;
        RECT 295.335 40.020 301.300 40.120 ;
        RECT 297.750 40.010 301.300 40.020 ;
        RECT 0.000 31.295 3.545 31.300 ;
        RECT 295.300 31.295 295.365 31.325 ;
        RECT 300.600 31.295 301.300 31.300 ;
        RECT 0.000 26.530 6.000 31.295 ;
        RECT 0.010 26.525 6.000 26.530 ;
        RECT 295.300 26.525 301.300 31.295 ;
        RECT 0.000 19.345 3.545 19.350 ;
        RECT 297.750 19.345 301.300 19.350 ;
        RECT 0.000 17.750 6.000 19.345 ;
        RECT 0.000 15.795 5.995 17.750 ;
        RECT 295.300 17.745 301.300 19.345 ;
        RECT 295.315 15.805 301.300 17.745 ;
        RECT 0.000 14.210 6.000 15.795 ;
        RECT 0.010 14.205 6.000 14.210 ;
        RECT 295.300 14.205 301.300 15.805 ;
        RECT 0.000 6.000 6.000 7.810 ;
        RECT 295.300 6.000 301.300 7.810 ;
        RECT 0.000 4.310 301.300 6.000 ;
        RECT 0.000 4.290 0.700 4.310 ;
        RECT 2.465 0.000 5.970 4.310 ;
        RECT 7.135 0.000 10.635 4.310 ;
        RECT 12.045 0.000 15.545 4.310 ;
        RECT 20.445 0.000 23.945 4.310 ;
        RECT 24.645 0.000 28.145 4.310 ;
        RECT 28.845 0.000 32.345 4.310 ;
        RECT 37.245 0.000 40.745 4.310 ;
        RECT 43.550 0.000 47.050 4.310 ;
        RECT 49.845 0.000 53.345 4.310 ;
        RECT 58.245 0.000 61.745 4.310 ;
        RECT 62.445 0.000 65.945 4.310 ;
        RECT 66.645 0.000 70.145 4.310 ;
        RECT 76.685 0.000 80.185 4.310 ;
        RECT 80.885 0.000 84.385 4.310 ;
        RECT 85.435 0.000 88.935 4.310 ;
        RECT 89.985 0.000 93.485 4.310 ;
        RECT 94.535 0.000 98.035 4.310 ;
        RECT 99.085 0.000 102.585 4.310 ;
        RECT 103.635 0.000 107.135 4.310 ;
        RECT 126.105 0.000 129.605 4.310 ;
        RECT 137.295 0.000 140.795 4.310 ;
        RECT 148.515 0.000 152.015 4.310 ;
        RECT 156.915 0.000 160.415 4.310 ;
        RECT 165.315 0.000 168.815 4.310 ;
        RECT 169.980 0.000 173.480 4.310 ;
        RECT 174.565 0.000 178.065 4.310 ;
        RECT 190.600 0.000 194.100 4.310 ;
        RECT 195.150 0.000 198.650 4.310 ;
        RECT 199.700 4.205 221.530 4.310 ;
        RECT 199.700 0.000 203.200 4.205 ;
        RECT 204.250 0.000 207.750 4.205 ;
        RECT 208.800 0.000 212.300 4.205 ;
        RECT 213.350 0.000 216.850 4.205 ;
        RECT 218.030 0.000 221.530 4.205 ;
        RECT 227.960 0.000 231.460 4.310 ;
        RECT 232.160 0.000 235.660 4.310 ;
        RECT 236.360 0.000 239.860 4.310 ;
        RECT 244.760 0.000 248.260 4.310 ;
        RECT 251.055 0.000 254.555 4.310 ;
        RECT 257.360 0.000 260.860 4.310 ;
        RECT 265.760 0.000 269.260 4.310 ;
        RECT 269.960 0.000 273.460 4.310 ;
        RECT 274.160 0.000 277.660 4.310 ;
        RECT 283.560 0.000 287.060 4.310 ;
        RECT 288.465 0.000 291.965 4.310 ;
        RECT 295.330 0.000 298.830 4.310 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.985 511.285 300.315 514.820 ;
        RECT 0.985 508.955 4.485 511.285 ;
        RECT 7.150 509.810 7.970 511.285 ;
        RECT 26.690 509.810 27.510 511.285 ;
        RECT 46.230 509.810 47.050 511.285 ;
        RECT 65.770 509.810 66.590 511.285 ;
        RECT 85.300 509.810 86.120 511.285 ;
        RECT 90.140 509.810 92.685 511.285 ;
        RECT 96.620 510.950 102.185 511.285 ;
        RECT 95.855 509.810 102.185 510.950 ;
        RECT 119.790 509.810 122.545 511.285 ;
        RECT 140.215 509.810 142.065 511.285 ;
        RECT 153.080 509.810 155.970 511.285 ;
        RECT 175.340 509.810 178.195 511.285 ;
        RECT 194.845 509.810 202.075 511.285 ;
        RECT 204.765 509.810 207.310 511.285 ;
        RECT 212.580 509.810 213.400 511.285 ;
        RECT 232.120 509.810 232.940 511.285 ;
        RECT 251.660 509.810 252.480 511.285 ;
        RECT 271.185 509.810 272.005 511.285 ;
        RECT 290.730 509.810 291.550 511.285 ;
        RECT 0.985 508.805 4.490 508.955 ;
        RECT 0.985 507.000 6.000 508.805 ;
        RECT 0.985 503.705 4.490 507.000 ;
        RECT 0.985 502.895 4.485 503.705 ;
        RECT 0.985 502.745 4.490 502.895 ;
        RECT 0.985 500.940 6.000 502.745 ;
        RECT 0.985 497.645 4.490 500.940 ;
        RECT 0.985 496.835 4.485 497.645 ;
        RECT 0.985 496.685 4.490 496.835 ;
        RECT 0.985 494.880 6.000 496.685 ;
        RECT 0.985 491.585 4.490 494.880 ;
        RECT 0.985 490.775 4.485 491.585 ;
        RECT 0.985 490.625 4.490 490.775 ;
        RECT 0.985 488.820 6.000 490.625 ;
        RECT 0.985 485.525 4.490 488.820 ;
        RECT 0.985 484.715 4.485 485.525 ;
        RECT 0.985 484.565 4.490 484.715 ;
        RECT 0.985 482.760 6.000 484.565 ;
        RECT 295.300 483.330 296.325 484.030 ;
        RECT 0.985 479.465 4.490 482.760 ;
        RECT 0.985 478.655 4.485 479.465 ;
        RECT 0.985 478.505 4.490 478.655 ;
        RECT 0.985 476.700 6.000 478.505 ;
        RECT 0.985 473.405 4.490 476.700 ;
        RECT 0.985 472.595 4.485 473.405 ;
        RECT 0.985 472.445 4.490 472.595 ;
        RECT 0.985 470.640 6.000 472.445 ;
        RECT 0.985 467.345 4.490 470.640 ;
        RECT 0.985 466.535 4.485 467.345 ;
        RECT 0.985 466.385 4.490 466.535 ;
        RECT 0.985 464.580 6.000 466.385 ;
        RECT 0.985 461.285 4.490 464.580 ;
        RECT 0.985 460.475 4.485 461.285 ;
        RECT 0.985 460.325 4.490 460.475 ;
        RECT 0.985 458.520 6.000 460.325 ;
        RECT 0.985 455.225 4.490 458.520 ;
        RECT 0.985 454.415 4.485 455.225 ;
        RECT 0.985 454.265 4.490 454.415 ;
        RECT 0.985 452.460 6.000 454.265 ;
        RECT 0.985 449.165 4.490 452.460 ;
        RECT 0.985 448.355 4.485 449.165 ;
        RECT 0.985 448.205 4.490 448.355 ;
        RECT 0.985 446.400 6.000 448.205 ;
        RECT 0.985 443.105 4.490 446.400 ;
        RECT 0.985 442.295 4.485 443.105 ;
        RECT 0.985 442.145 4.490 442.295 ;
        RECT 0.985 440.340 6.000 442.145 ;
        RECT 0.985 437.045 4.490 440.340 ;
        RECT 0.985 436.235 4.485 437.045 ;
        RECT 0.985 436.085 4.490 436.235 ;
        RECT 0.985 434.280 6.000 436.085 ;
        RECT 0.985 430.985 4.490 434.280 ;
        RECT 0.985 430.175 4.485 430.985 ;
        RECT 0.985 430.025 4.490 430.175 ;
        RECT 0.985 428.220 6.000 430.025 ;
        RECT 0.985 424.925 4.490 428.220 ;
        RECT 0.985 424.115 4.485 424.925 ;
        RECT 0.985 423.965 4.490 424.115 ;
        RECT 0.985 422.160 6.000 423.965 ;
        RECT 0.985 418.865 4.490 422.160 ;
        RECT 0.985 418.055 4.485 418.865 ;
        RECT 0.985 417.905 4.490 418.055 ;
        RECT 0.985 416.100 6.000 417.905 ;
        RECT 0.985 412.805 4.490 416.100 ;
        RECT 0.985 411.995 4.485 412.805 ;
        RECT 0.985 411.845 4.490 411.995 ;
        RECT 0.985 410.040 6.000 411.845 ;
        RECT 0.985 406.745 4.490 410.040 ;
        RECT 0.985 405.935 4.485 406.745 ;
        RECT 0.985 405.785 4.490 405.935 ;
        RECT 0.985 403.980 6.000 405.785 ;
        RECT 0.985 400.685 4.490 403.980 ;
        RECT 0.985 399.875 4.485 400.685 ;
        RECT 0.985 399.725 4.490 399.875 ;
        RECT 0.985 397.920 6.000 399.725 ;
        RECT 0.985 394.625 4.490 397.920 ;
        RECT 0.985 393.815 4.485 394.625 ;
        RECT 0.985 393.665 4.490 393.815 ;
        RECT 0.985 391.860 6.000 393.665 ;
        RECT 0.985 388.565 4.490 391.860 ;
        RECT 0.985 387.755 4.485 388.565 ;
        RECT 0.985 387.605 4.490 387.755 ;
        RECT 0.985 385.800 6.000 387.605 ;
        RECT 0.985 382.505 4.490 385.800 ;
        RECT 0.985 381.695 4.485 382.505 ;
        RECT 0.985 381.545 4.490 381.695 ;
        RECT 0.985 379.740 6.000 381.545 ;
        RECT 0.985 376.445 4.490 379.740 ;
        RECT 0.985 375.635 4.485 376.445 ;
        RECT 0.985 375.485 4.490 375.635 ;
        RECT 0.985 373.680 6.000 375.485 ;
        RECT 0.985 370.385 4.490 373.680 ;
        RECT 0.985 369.575 4.485 370.385 ;
        RECT 0.985 369.425 4.490 369.575 ;
        RECT 0.985 367.620 6.000 369.425 ;
        RECT 0.985 364.325 4.490 367.620 ;
        RECT 0.985 363.515 4.485 364.325 ;
        RECT 0.985 363.365 4.490 363.515 ;
        RECT 0.985 361.560 6.000 363.365 ;
        RECT 0.985 358.265 4.490 361.560 ;
        RECT 0.985 357.455 4.485 358.265 ;
        RECT 0.985 357.305 4.490 357.455 ;
        RECT 0.985 355.500 6.000 357.305 ;
        RECT 0.985 352.205 4.490 355.500 ;
        RECT 0.985 351.395 4.485 352.205 ;
        RECT 0.985 351.245 4.490 351.395 ;
        RECT 0.985 349.440 6.000 351.245 ;
        RECT 0.985 346.145 4.490 349.440 ;
        RECT 0.985 345.335 4.485 346.145 ;
        RECT 0.985 345.185 4.490 345.335 ;
        RECT 0.985 343.380 6.000 345.185 ;
        RECT 0.985 340.085 4.490 343.380 ;
        RECT 0.985 339.275 4.485 340.085 ;
        RECT 0.985 339.125 4.490 339.275 ;
        RECT 0.985 337.320 6.000 339.125 ;
        RECT 0.985 334.025 4.490 337.320 ;
        RECT 0.985 333.215 4.485 334.025 ;
        RECT 0.985 333.065 4.490 333.215 ;
        RECT 0.985 331.260 6.000 333.065 ;
        RECT 0.985 327.965 4.490 331.260 ;
        RECT 0.985 327.155 4.485 327.965 ;
        RECT 0.985 327.005 4.490 327.155 ;
        RECT 0.985 325.200 6.000 327.005 ;
        RECT 0.985 321.905 4.490 325.200 ;
        RECT 0.985 321.095 4.485 321.905 ;
        RECT 0.985 320.945 4.490 321.095 ;
        RECT 0.985 319.140 6.000 320.945 ;
        RECT 0.985 315.845 4.490 319.140 ;
        RECT 0.985 315.035 4.485 315.845 ;
        RECT 0.985 314.885 4.490 315.035 ;
        RECT 0.985 313.080 6.000 314.885 ;
        RECT 0.985 309.785 4.490 313.080 ;
        RECT 0.985 308.975 4.485 309.785 ;
        RECT 0.985 308.825 4.490 308.975 ;
        RECT 0.985 307.020 6.000 308.825 ;
        RECT 0.985 303.725 4.490 307.020 ;
        RECT 0.985 302.915 4.485 303.725 ;
        RECT 0.985 302.765 4.490 302.915 ;
        RECT 0.985 300.960 6.000 302.765 ;
        RECT 0.985 297.665 4.490 300.960 ;
        RECT 0.985 296.855 4.485 297.665 ;
        RECT 0.985 296.705 4.490 296.855 ;
        RECT 0.985 294.900 6.000 296.705 ;
        RECT 0.985 291.605 4.490 294.900 ;
        RECT 0.985 290.795 4.485 291.605 ;
        RECT 0.985 290.645 4.490 290.795 ;
        RECT 0.985 288.840 6.000 290.645 ;
        RECT 0.985 285.545 4.490 288.840 ;
        RECT 0.985 284.735 4.485 285.545 ;
        RECT 0.985 284.585 4.490 284.735 ;
        RECT 0.985 282.780 6.000 284.585 ;
        RECT 0.985 279.485 4.490 282.780 ;
        RECT 0.985 278.675 4.485 279.485 ;
        RECT 0.985 278.525 4.490 278.675 ;
        RECT 0.985 276.720 6.000 278.525 ;
        RECT 0.985 273.425 4.490 276.720 ;
        RECT 0.985 272.615 4.485 273.425 ;
        RECT 0.985 272.465 4.490 272.615 ;
        RECT 0.985 270.660 6.000 272.465 ;
        RECT 0.985 267.365 4.490 270.660 ;
        RECT 0.985 266.555 4.485 267.365 ;
        RECT 0.985 266.405 4.490 266.555 ;
        RECT 0.985 264.600 6.000 266.405 ;
        RECT 0.985 261.305 4.490 264.600 ;
        RECT 0.985 260.495 4.485 261.305 ;
        RECT 0.985 260.345 4.490 260.495 ;
        RECT 0.985 258.540 6.000 260.345 ;
        RECT 0.985 255.245 4.490 258.540 ;
        RECT 0.985 254.435 4.485 255.245 ;
        RECT 0.985 254.285 4.490 254.435 ;
        RECT 0.985 252.480 6.000 254.285 ;
        RECT 0.985 249.185 4.490 252.480 ;
        RECT 0.985 248.375 4.485 249.185 ;
        RECT 0.985 248.225 4.490 248.375 ;
        RECT 0.985 246.420 6.000 248.225 ;
        RECT 0.985 243.125 4.490 246.420 ;
        RECT 0.985 242.315 4.485 243.125 ;
        RECT 0.985 242.165 4.490 242.315 ;
        RECT 0.985 240.360 6.000 242.165 ;
        RECT 0.985 237.065 4.490 240.360 ;
        RECT 0.985 236.255 4.485 237.065 ;
        RECT 0.985 236.105 4.490 236.255 ;
        RECT 0.985 234.300 6.000 236.105 ;
        RECT 0.985 231.005 4.490 234.300 ;
        RECT 0.985 230.195 4.485 231.005 ;
        RECT 0.985 230.045 4.490 230.195 ;
        RECT 0.985 228.240 6.000 230.045 ;
        RECT 0.985 224.945 4.490 228.240 ;
        RECT 0.985 224.135 4.485 224.945 ;
        RECT 0.985 223.985 4.490 224.135 ;
        RECT 0.985 222.180 6.000 223.985 ;
        RECT 0.985 218.885 4.490 222.180 ;
        RECT 0.985 218.075 4.485 218.885 ;
        RECT 0.985 217.925 4.490 218.075 ;
        RECT 0.985 216.120 6.000 217.925 ;
        RECT 0.985 212.825 4.490 216.120 ;
        RECT 0.985 212.015 4.485 212.825 ;
        RECT 0.985 211.865 4.490 212.015 ;
        RECT 0.985 210.060 6.000 211.865 ;
        RECT 0.985 206.765 4.490 210.060 ;
        RECT 0.985 205.955 4.485 206.765 ;
        RECT 0.985 205.805 4.490 205.955 ;
        RECT 0.985 204.000 6.000 205.805 ;
        RECT 0.985 200.705 4.490 204.000 ;
        RECT 0.985 199.895 4.485 200.705 ;
        RECT 0.985 199.745 4.490 199.895 ;
        RECT 0.985 197.940 6.000 199.745 ;
        RECT 0.985 194.645 4.490 197.940 ;
        RECT 0.985 193.835 4.485 194.645 ;
        RECT 0.985 193.685 4.490 193.835 ;
        RECT 0.985 191.880 6.000 193.685 ;
        RECT 0.985 188.585 4.490 191.880 ;
        RECT 0.985 187.775 4.485 188.585 ;
        RECT 0.985 187.625 4.490 187.775 ;
        RECT 0.985 185.820 6.000 187.625 ;
        RECT 0.985 182.525 4.490 185.820 ;
        RECT 0.985 181.715 4.485 182.525 ;
        RECT 0.985 181.565 4.490 181.715 ;
        RECT 0.985 179.760 6.000 181.565 ;
        RECT 0.985 176.465 4.490 179.760 ;
        RECT 0.985 175.655 4.485 176.465 ;
        RECT 0.985 175.505 4.490 175.655 ;
        RECT 0.985 173.700 6.000 175.505 ;
        RECT 0.985 170.405 4.490 173.700 ;
        RECT 0.985 169.595 4.485 170.405 ;
        RECT 0.985 169.445 4.490 169.595 ;
        RECT 0.985 167.640 6.000 169.445 ;
        RECT 0.985 164.345 4.490 167.640 ;
        RECT 0.985 163.535 4.485 164.345 ;
        RECT 0.985 163.385 4.490 163.535 ;
        RECT 0.985 161.580 6.000 163.385 ;
        RECT 0.985 158.285 4.490 161.580 ;
        RECT 0.985 157.475 4.485 158.285 ;
        RECT 0.985 157.325 4.490 157.475 ;
        RECT 0.985 155.520 6.000 157.325 ;
        RECT 0.985 152.225 4.490 155.520 ;
        RECT 0.985 151.415 4.485 152.225 ;
        RECT 0.985 151.265 4.490 151.415 ;
        RECT 0.985 149.460 6.000 151.265 ;
        RECT 0.985 146.165 4.490 149.460 ;
        RECT 0.985 145.355 4.485 146.165 ;
        RECT 0.985 145.205 4.490 145.355 ;
        RECT 0.985 143.400 6.000 145.205 ;
        RECT 0.985 140.105 4.490 143.400 ;
        RECT 0.985 139.295 4.485 140.105 ;
        RECT 0.985 139.145 4.490 139.295 ;
        RECT 0.985 137.340 6.000 139.145 ;
        RECT 0.985 134.045 4.490 137.340 ;
        RECT 0.985 133.235 4.485 134.045 ;
        RECT 0.985 133.085 4.490 133.235 ;
        RECT 0.985 131.280 6.000 133.085 ;
        RECT 0.985 127.985 4.490 131.280 ;
        RECT 0.985 127.175 4.485 127.985 ;
        RECT 0.985 127.025 4.490 127.175 ;
        RECT 0.985 125.220 6.000 127.025 ;
        RECT 0.985 121.925 4.490 125.220 ;
        RECT 0.985 121.115 4.485 121.925 ;
        RECT 0.985 120.965 4.490 121.115 ;
        RECT 0.985 119.160 6.000 120.965 ;
        RECT 0.985 115.865 4.490 119.160 ;
        RECT 0.985 87.265 4.485 115.865 ;
        RECT 296.815 114.965 300.315 511.285 ;
        RECT 295.300 114.355 300.315 114.965 ;
        RECT 296.815 112.405 300.315 114.355 ;
        RECT 295.300 111.810 300.315 112.405 ;
        RECT 296.815 87.265 300.315 111.810 ;
        RECT 0.985 86.795 6.000 87.265 ;
        RECT 295.300 86.795 300.315 87.265 ;
        RECT 0.985 72.515 4.485 86.795 ;
        RECT 296.815 72.515 300.315 86.795 ;
        RECT 0.985 71.835 6.000 72.515 ;
        RECT 295.300 71.835 300.315 72.515 ;
        RECT 0.985 4.485 4.485 71.835 ;
        RECT 95.850 4.485 202.075 6.000 ;
        RECT 296.815 4.485 300.315 71.835 ;
        RECT 0.985 4.480 202.505 4.485 ;
        RECT 204.680 4.480 300.315 4.485 ;
        RECT 0.985 0.985 300.315 4.480 ;
        RECT 87.030 0.980 87.730 0.985 ;
        RECT 90.590 0.980 91.290 0.985 ;
      LAYER Metal2 ;
        RECT 0.985 513.680 300.315 514.820 ;
        RECT 0.995 506.690 2.125 509.120 ;
        RECT 299.120 506.675 300.800 509.105 ;
        RECT 0.995 500.630 2.125 503.060 ;
        RECT 299.120 500.615 300.800 503.045 ;
        RECT 0.995 494.570 2.125 497.000 ;
        RECT 299.120 494.555 300.800 496.985 ;
        RECT 0.995 488.510 2.125 490.940 ;
        RECT 299.120 488.495 300.800 490.925 ;
        RECT 0.995 482.450 2.125 484.880 ;
        RECT 299.120 482.435 300.800 484.865 ;
        RECT 0.995 476.390 2.125 478.820 ;
        RECT 299.120 476.375 300.800 478.805 ;
        RECT 0.995 470.330 2.125 472.760 ;
        RECT 299.120 470.315 300.800 472.745 ;
        RECT 0.995 464.270 2.125 466.700 ;
        RECT 299.120 464.255 300.800 466.685 ;
        RECT 0.995 458.210 2.125 460.640 ;
        RECT 299.120 458.195 300.800 460.625 ;
        RECT 0.995 452.150 2.125 454.580 ;
        RECT 299.120 452.135 300.800 454.565 ;
        RECT 0.995 446.090 2.125 448.520 ;
        RECT 299.120 446.075 300.800 448.505 ;
        RECT 0.995 440.030 2.125 442.460 ;
        RECT 299.120 440.015 300.800 442.445 ;
        RECT 0.995 433.970 2.125 436.400 ;
        RECT 299.120 433.955 300.800 436.385 ;
        RECT 0.995 427.910 2.125 430.340 ;
        RECT 299.120 427.895 300.800 430.325 ;
        RECT 0.995 421.850 2.125 424.280 ;
        RECT 299.120 421.835 300.800 424.265 ;
        RECT 0.995 415.790 2.125 418.220 ;
        RECT 299.120 415.775 300.800 418.205 ;
        RECT 0.995 409.730 2.125 412.160 ;
        RECT 299.120 409.715 300.800 412.145 ;
        RECT 0.995 403.670 2.125 406.100 ;
        RECT 299.120 403.655 300.800 406.085 ;
        RECT 0.995 397.610 2.125 400.040 ;
        RECT 299.120 397.595 300.800 400.025 ;
        RECT 0.995 391.550 2.125 393.980 ;
        RECT 299.120 391.535 300.800 393.965 ;
        RECT 0.995 385.490 2.125 387.920 ;
        RECT 299.120 385.475 300.800 387.905 ;
        RECT 0.995 379.430 2.125 381.860 ;
        RECT 299.120 379.415 300.800 381.845 ;
        RECT 0.995 373.370 2.125 375.800 ;
        RECT 299.120 373.355 300.800 375.785 ;
        RECT 0.995 367.310 2.125 369.740 ;
        RECT 299.120 367.295 300.800 369.725 ;
        RECT 0.995 361.250 2.125 363.680 ;
        RECT 299.120 361.235 300.800 363.665 ;
        RECT 0.995 355.190 2.125 357.620 ;
        RECT 299.120 355.175 300.800 357.605 ;
        RECT 0.995 349.130 2.125 351.560 ;
        RECT 299.120 349.115 300.800 351.545 ;
        RECT 0.995 343.070 2.125 345.500 ;
        RECT 299.120 343.055 300.800 345.485 ;
        RECT 0.995 337.010 2.125 339.440 ;
        RECT 299.120 336.995 300.800 339.425 ;
        RECT 0.995 330.950 2.125 333.380 ;
        RECT 299.120 330.935 300.800 333.365 ;
        RECT 0.995 324.890 2.125 327.320 ;
        RECT 299.120 324.875 300.800 327.305 ;
        RECT 0.995 318.830 2.125 321.260 ;
        RECT 299.120 318.815 300.800 321.245 ;
        RECT 0.995 312.770 2.125 315.200 ;
        RECT 299.120 312.755 300.800 315.185 ;
        RECT 0.995 306.710 2.125 309.140 ;
        RECT 299.120 306.695 300.800 309.125 ;
        RECT 0.995 300.650 2.125 303.080 ;
        RECT 299.120 300.635 300.800 303.065 ;
        RECT 0.995 294.590 2.125 297.020 ;
        RECT 299.120 294.575 300.800 297.005 ;
        RECT 0.995 288.530 2.125 290.960 ;
        RECT 299.120 288.515 300.800 290.945 ;
        RECT 0.995 282.470 2.125 284.900 ;
        RECT 299.120 282.455 300.800 284.885 ;
        RECT 0.995 276.410 2.125 278.840 ;
        RECT 299.120 276.395 300.800 278.825 ;
        RECT 0.995 270.350 2.125 272.780 ;
        RECT 299.120 270.335 300.800 272.765 ;
        RECT 0.995 264.290 2.125 266.720 ;
        RECT 299.120 264.275 300.800 266.705 ;
        RECT 0.995 258.230 2.125 260.660 ;
        RECT 299.120 258.215 300.800 260.645 ;
        RECT 0.995 252.170 2.125 254.600 ;
        RECT 299.120 252.155 300.800 254.585 ;
        RECT 0.995 246.110 2.125 248.540 ;
        RECT 299.120 246.095 300.800 248.525 ;
        RECT 0.995 240.050 2.125 242.480 ;
        RECT 299.120 240.035 300.800 242.465 ;
        RECT 0.995 233.990 2.125 236.420 ;
        RECT 299.120 233.975 300.800 236.405 ;
        RECT 0.995 227.930 2.125 230.360 ;
        RECT 299.120 227.915 300.800 230.345 ;
        RECT 0.995 221.870 2.125 224.300 ;
        RECT 299.120 221.855 300.800 224.285 ;
        RECT 0.995 215.810 2.125 218.240 ;
        RECT 299.120 215.795 300.800 218.225 ;
        RECT 0.995 209.750 2.125 212.180 ;
        RECT 299.120 209.735 300.800 212.165 ;
        RECT 0.995 203.690 2.125 206.120 ;
        RECT 299.120 203.675 300.800 206.105 ;
        RECT 0.995 197.630 2.125 200.060 ;
        RECT 299.120 197.615 300.800 200.045 ;
        RECT 0.995 191.570 2.125 194.000 ;
        RECT 299.120 191.555 300.800 193.985 ;
        RECT 0.995 185.510 2.125 187.940 ;
        RECT 299.120 185.495 300.800 187.925 ;
        RECT 0.995 179.450 2.125 181.880 ;
        RECT 299.120 179.435 300.800 181.865 ;
        RECT 0.995 173.390 2.125 175.820 ;
        RECT 299.120 173.375 300.800 175.805 ;
        RECT 0.995 167.330 2.125 169.760 ;
        RECT 299.120 167.315 300.800 169.745 ;
        RECT 0.995 161.270 2.125 163.700 ;
        RECT 299.120 161.255 300.800 163.685 ;
        RECT 0.995 155.210 2.125 157.640 ;
        RECT 299.120 155.195 300.800 157.625 ;
        RECT 0.995 149.150 2.125 151.580 ;
        RECT 299.120 149.135 300.800 151.565 ;
        RECT 0.995 143.090 2.125 145.520 ;
        RECT 299.120 143.075 300.800 145.505 ;
        RECT 0.995 137.030 2.125 139.460 ;
        RECT 299.120 137.015 300.800 139.445 ;
        RECT 0.995 130.970 2.125 133.400 ;
        RECT 299.120 130.955 300.800 133.385 ;
        RECT 0.995 124.910 2.125 127.340 ;
        RECT 299.120 124.895 300.800 127.325 ;
        RECT 0.995 118.850 2.125 121.280 ;
        RECT 299.120 118.835 300.800 121.265 ;
        RECT 0.995 111.495 2.125 113.925 ;
        RECT 299.185 111.495 300.315 113.925 ;
        RECT 0.995 83.455 2.125 92.695 ;
        RECT 299.185 83.455 300.315 92.695 ;
        RECT 0.995 69.460 2.125 72.760 ;
        RECT 299.185 69.460 300.315 72.760 ;
        RECT 0.995 48.095 2.125 57.145 ;
        RECT 299.185 48.095 300.315 57.145 ;
        RECT 0.995 33.790 2.125 37.960 ;
        RECT 299.185 33.790 300.315 37.960 ;
        RECT 0.995 19.880 2.125 26.220 ;
        RECT 299.185 19.880 300.315 26.220 ;
        RECT 0.995 8.890 2.125 13.060 ;
        RECT 299.185 8.890 300.315 13.060 ;
        RECT 16.245 0.985 19.745 4.485 ;
        RECT 25.040 0.985 25.820 6.000 ;
        RECT 28.600 0.985 29.385 6.000 ;
        RECT 33.045 0.985 36.545 4.485 ;
        RECT 54.045 0.985 57.545 4.485 ;
        RECT 63.850 0.985 64.630 6.000 ;
        RECT 67.410 0.985 68.195 6.000 ;
        RECT 70.845 0.985 74.345 4.485 ;
        RECT 87.000 0.975 87.775 6.000 ;
        RECT 90.555 0.975 91.335 6.000 ;
        RECT 109.630 0.985 113.130 4.485 ;
        RECT 115.575 0.985 119.075 4.485 ;
        RECT 121.905 0.985 125.405 4.485 ;
        RECT 129.495 4.310 130.275 6.000 ;
        RECT 133.055 4.485 133.840 6.000 ;
        RECT 135.865 4.485 136.645 6.000 ;
        RECT 133.055 4.310 136.645 4.485 ;
        RECT 139.425 4.310 140.210 6.000 ;
        RECT 133.095 0.985 136.595 4.310 ;
        RECT 144.315 0.985 147.815 4.485 ;
        RECT 152.715 0.985 156.215 4.485 ;
        RECT 161.115 0.985 164.615 4.485 ;
        RECT 179.315 0.985 182.815 4.485 ;
        RECT 183.670 0.985 187.170 4.485 ;
        RECT 206.100 1.005 206.875 6.000 ;
        RECT 209.655 1.005 210.435 6.000 ;
        RECT 223.760 0.985 227.260 4.485 ;
        RECT 230.315 0.985 231.095 6.000 ;
        RECT 233.875 0.985 234.660 6.000 ;
        RECT 240.560 0.985 244.060 4.485 ;
        RECT 261.560 0.985 265.060 4.485 ;
        RECT 269.465 0.965 270.245 6.000 ;
        RECT 273.025 0.965 273.810 6.000 ;
        RECT 278.360 0.985 281.860 4.485 ;
      LAYER Metal3 ;
        RECT 9.370 513.675 12.870 515.810 ;
        RECT 18.760 513.680 22.260 515.810 ;
        RECT 28.910 513.675 32.410 515.810 ;
        RECT 37.660 513.680 41.160 515.810 ;
        RECT 48.450 513.675 51.950 515.810 ;
        RECT 56.560 513.680 60.060 515.810 ;
        RECT 67.990 513.675 71.490 515.810 ;
        RECT 80.400 513.675 83.900 515.810 ;
        RECT 88.805 513.680 92.305 515.810 ;
        RECT 98.320 513.680 101.820 515.810 ;
        RECT 103.205 513.680 106.705 515.810 ;
        RECT 114.085 513.680 117.585 515.810 ;
        RECT 119.835 513.680 123.335 515.810 ;
        RECT 130.070 513.680 133.570 515.810 ;
        RECT 140.340 513.680 143.840 515.810 ;
        RECT 149.255 513.680 152.755 515.810 ;
        RECT 153.745 513.680 157.245 515.810 ;
        RECT 166.375 513.680 169.875 515.810 ;
        RECT 177.380 513.680 180.880 515.810 ;
        RECT 196.715 513.680 200.215 515.810 ;
        RECT 205.520 513.680 209.020 515.810 ;
        RECT 214.800 513.675 218.300 515.810 ;
        RECT 226.275 513.680 229.775 515.810 ;
        RECT 234.340 513.675 237.840 515.810 ;
        RECT 245.175 513.680 248.675 515.810 ;
        RECT 253.880 513.675 257.380 515.810 ;
        RECT 264.075 513.680 267.575 515.810 ;
        RECT 273.405 513.675 276.905 515.810 ;
        RECT 285.830 513.675 289.330 515.810 ;
        RECT 0.000 508.430 3.555 509.130 ;
        RECT 297.755 509.010 301.300 509.115 ;
        RECT 297.750 508.615 301.300 509.010 ;
        RECT 0.000 507.380 6.000 508.430 ;
        RECT 295.300 507.565 301.300 508.615 ;
        RECT 0.000 506.680 3.555 507.380 ;
        RECT 297.750 506.565 301.300 507.565 ;
        RECT 0.000 502.370 3.555 503.070 ;
        RECT 297.755 502.950 301.300 503.055 ;
        RECT 297.750 502.555 301.300 502.950 ;
        RECT 0.000 501.320 6.000 502.370 ;
        RECT 295.300 501.505 301.300 502.555 ;
        RECT 0.000 500.620 3.555 501.320 ;
        RECT 297.750 500.505 301.300 501.505 ;
        RECT 0.000 496.310 3.555 497.010 ;
        RECT 297.755 496.890 301.300 496.995 ;
        RECT 297.750 496.495 301.300 496.890 ;
        RECT 0.000 495.260 6.000 496.310 ;
        RECT 295.300 495.445 301.300 496.495 ;
        RECT 0.000 494.560 3.555 495.260 ;
        RECT 297.750 494.445 301.300 495.445 ;
        RECT 0.000 490.250 3.555 490.950 ;
        RECT 297.755 490.830 301.300 490.935 ;
        RECT 297.750 490.435 301.300 490.830 ;
        RECT 0.000 489.200 6.000 490.250 ;
        RECT 295.300 489.385 301.300 490.435 ;
        RECT 0.000 488.500 3.555 489.200 ;
        RECT 297.750 488.385 301.300 489.385 ;
        RECT 0.000 484.190 3.555 484.890 ;
        RECT 297.755 484.770 301.300 484.875 ;
        RECT 297.750 484.375 301.300 484.770 ;
        RECT 0.000 483.140 6.000 484.190 ;
        RECT 295.300 483.325 301.300 484.375 ;
        RECT 0.000 482.440 3.555 483.140 ;
        RECT 297.750 482.325 301.300 483.325 ;
        RECT 0.000 478.130 3.555 478.830 ;
        RECT 297.755 478.710 301.300 478.815 ;
        RECT 297.750 478.315 301.300 478.710 ;
        RECT 0.000 477.080 6.000 478.130 ;
        RECT 295.300 477.265 301.300 478.315 ;
        RECT 0.000 476.380 3.555 477.080 ;
        RECT 297.750 476.265 301.300 477.265 ;
        RECT 0.000 472.070 3.555 472.770 ;
        RECT 297.755 472.650 301.300 472.755 ;
        RECT 297.750 472.255 301.300 472.650 ;
        RECT 0.000 471.020 6.000 472.070 ;
        RECT 295.300 471.205 301.300 472.255 ;
        RECT 0.000 470.320 3.555 471.020 ;
        RECT 297.750 470.205 301.300 471.205 ;
        RECT 0.000 466.010 3.555 466.710 ;
        RECT 297.755 466.590 301.300 466.695 ;
        RECT 297.750 466.195 301.300 466.590 ;
        RECT 0.000 464.960 6.000 466.010 ;
        RECT 295.300 465.145 301.300 466.195 ;
        RECT 0.000 464.260 3.555 464.960 ;
        RECT 297.750 464.145 301.300 465.145 ;
        RECT 0.000 459.950 3.555 460.650 ;
        RECT 297.755 460.530 301.300 460.635 ;
        RECT 297.750 460.135 301.300 460.530 ;
        RECT 0.000 458.900 6.000 459.950 ;
        RECT 295.300 459.085 301.300 460.135 ;
        RECT 0.000 458.200 3.555 458.900 ;
        RECT 297.750 458.085 301.300 459.085 ;
        RECT 0.000 453.890 3.555 454.590 ;
        RECT 297.755 454.470 301.300 454.575 ;
        RECT 297.750 454.075 301.300 454.470 ;
        RECT 0.000 452.840 6.000 453.890 ;
        RECT 295.300 453.025 301.300 454.075 ;
        RECT 0.000 452.140 3.555 452.840 ;
        RECT 297.750 452.025 301.300 453.025 ;
        RECT 0.000 447.830 3.555 448.530 ;
        RECT 297.755 448.410 301.300 448.515 ;
        RECT 297.750 448.015 301.300 448.410 ;
        RECT 0.000 446.780 6.000 447.830 ;
        RECT 295.300 446.965 301.300 448.015 ;
        RECT 0.000 446.080 3.555 446.780 ;
        RECT 297.750 445.965 301.300 446.965 ;
        RECT 0.000 441.770 3.555 442.470 ;
        RECT 297.755 442.350 301.300 442.455 ;
        RECT 297.750 441.955 301.300 442.350 ;
        RECT 0.000 440.720 6.000 441.770 ;
        RECT 295.300 440.905 301.300 441.955 ;
        RECT 0.000 440.020 3.555 440.720 ;
        RECT 297.750 439.905 301.300 440.905 ;
        RECT 0.000 435.710 3.555 436.410 ;
        RECT 297.755 436.290 301.300 436.395 ;
        RECT 297.750 435.895 301.300 436.290 ;
        RECT 0.000 434.660 6.000 435.710 ;
        RECT 295.300 434.845 301.300 435.895 ;
        RECT 0.000 433.960 3.555 434.660 ;
        RECT 297.750 433.845 301.300 434.845 ;
        RECT 0.000 429.650 3.555 430.350 ;
        RECT 297.755 430.230 301.300 430.335 ;
        RECT 297.750 429.835 301.300 430.230 ;
        RECT 0.000 428.600 6.000 429.650 ;
        RECT 295.300 428.785 301.300 429.835 ;
        RECT 0.000 427.900 3.555 428.600 ;
        RECT 297.750 427.785 301.300 428.785 ;
        RECT 0.000 423.590 3.555 424.290 ;
        RECT 297.755 424.170 301.300 424.275 ;
        RECT 297.750 423.775 301.300 424.170 ;
        RECT 0.000 422.540 6.000 423.590 ;
        RECT 295.300 422.725 301.300 423.775 ;
        RECT 0.000 421.840 3.555 422.540 ;
        RECT 297.750 421.725 301.300 422.725 ;
        RECT 0.000 417.530 3.555 418.230 ;
        RECT 297.755 418.110 301.300 418.215 ;
        RECT 297.750 417.715 301.300 418.110 ;
        RECT 0.000 416.480 6.000 417.530 ;
        RECT 295.300 416.665 301.300 417.715 ;
        RECT 0.000 415.780 3.555 416.480 ;
        RECT 297.750 415.665 301.300 416.665 ;
        RECT 0.000 411.470 3.555 412.170 ;
        RECT 297.755 412.050 301.300 412.155 ;
        RECT 297.750 411.655 301.300 412.050 ;
        RECT 0.000 410.420 6.000 411.470 ;
        RECT 295.300 410.605 301.300 411.655 ;
        RECT 0.000 409.720 3.555 410.420 ;
        RECT 297.750 409.605 301.300 410.605 ;
        RECT 0.000 405.410 3.555 406.110 ;
        RECT 297.755 405.990 301.300 406.095 ;
        RECT 297.750 405.595 301.300 405.990 ;
        RECT 0.000 404.360 6.000 405.410 ;
        RECT 295.300 404.545 301.300 405.595 ;
        RECT 0.000 403.660 3.555 404.360 ;
        RECT 297.750 403.545 301.300 404.545 ;
        RECT 0.000 399.350 3.555 400.050 ;
        RECT 297.755 399.930 301.300 400.035 ;
        RECT 297.750 399.535 301.300 399.930 ;
        RECT 0.000 398.300 6.000 399.350 ;
        RECT 295.300 398.485 301.300 399.535 ;
        RECT 0.000 397.600 3.555 398.300 ;
        RECT 297.750 397.485 301.300 398.485 ;
        RECT 0.000 393.290 3.555 393.990 ;
        RECT 297.755 393.870 301.300 393.975 ;
        RECT 297.750 393.475 301.300 393.870 ;
        RECT 0.000 392.240 6.000 393.290 ;
        RECT 295.300 392.425 301.300 393.475 ;
        RECT 0.000 391.540 3.555 392.240 ;
        RECT 297.750 391.425 301.300 392.425 ;
        RECT 0.000 387.230 3.555 387.930 ;
        RECT 297.755 387.810 301.300 387.915 ;
        RECT 297.750 387.415 301.300 387.810 ;
        RECT 0.000 386.180 6.000 387.230 ;
        RECT 295.300 386.365 301.300 387.415 ;
        RECT 0.000 385.480 3.555 386.180 ;
        RECT 297.750 385.365 301.300 386.365 ;
        RECT 0.000 381.170 3.555 381.870 ;
        RECT 297.755 381.750 301.300 381.855 ;
        RECT 297.750 381.355 301.300 381.750 ;
        RECT 0.000 380.120 6.000 381.170 ;
        RECT 295.300 380.305 301.300 381.355 ;
        RECT 0.000 379.420 3.555 380.120 ;
        RECT 297.750 379.305 301.300 380.305 ;
        RECT 0.000 375.110 3.555 375.810 ;
        RECT 297.755 375.690 301.300 375.795 ;
        RECT 297.750 375.295 301.300 375.690 ;
        RECT 0.000 374.060 6.000 375.110 ;
        RECT 295.300 374.245 301.300 375.295 ;
        RECT 0.000 373.360 3.555 374.060 ;
        RECT 297.750 373.245 301.300 374.245 ;
        RECT 0.000 369.050 3.555 369.750 ;
        RECT 297.755 369.630 301.300 369.735 ;
        RECT 297.750 369.235 301.300 369.630 ;
        RECT 0.000 368.000 6.000 369.050 ;
        RECT 295.300 368.185 301.300 369.235 ;
        RECT 0.000 367.300 3.555 368.000 ;
        RECT 297.750 367.185 301.300 368.185 ;
        RECT 0.000 362.990 3.555 363.690 ;
        RECT 297.755 363.570 301.300 363.675 ;
        RECT 297.750 363.175 301.300 363.570 ;
        RECT 0.000 361.940 6.000 362.990 ;
        RECT 295.300 362.125 301.300 363.175 ;
        RECT 0.000 361.240 3.555 361.940 ;
        RECT 297.750 361.125 301.300 362.125 ;
        RECT 0.000 356.930 3.555 357.630 ;
        RECT 297.755 357.510 301.300 357.615 ;
        RECT 297.750 357.115 301.300 357.510 ;
        RECT 0.000 355.880 6.000 356.930 ;
        RECT 295.300 356.065 301.300 357.115 ;
        RECT 0.000 355.180 3.555 355.880 ;
        RECT 297.750 355.065 301.300 356.065 ;
        RECT 0.000 350.870 3.555 351.570 ;
        RECT 297.755 351.450 301.300 351.555 ;
        RECT 297.750 351.055 301.300 351.450 ;
        RECT 0.000 349.820 6.000 350.870 ;
        RECT 295.300 350.005 301.300 351.055 ;
        RECT 0.000 349.120 3.555 349.820 ;
        RECT 297.750 349.005 301.300 350.005 ;
        RECT 0.000 344.810 3.555 345.510 ;
        RECT 297.755 345.390 301.300 345.495 ;
        RECT 297.750 344.995 301.300 345.390 ;
        RECT 0.000 343.760 6.000 344.810 ;
        RECT 295.300 343.945 301.300 344.995 ;
        RECT 0.000 343.060 3.555 343.760 ;
        RECT 297.750 342.945 301.300 343.945 ;
        RECT 0.000 338.750 3.555 339.450 ;
        RECT 297.755 339.330 301.300 339.435 ;
        RECT 297.750 338.935 301.300 339.330 ;
        RECT 0.000 337.700 6.000 338.750 ;
        RECT 295.300 337.885 301.300 338.935 ;
        RECT 0.000 337.000 3.555 337.700 ;
        RECT 297.750 336.885 301.300 337.885 ;
        RECT 0.000 332.690 3.555 333.390 ;
        RECT 297.755 333.270 301.300 333.375 ;
        RECT 297.750 332.875 301.300 333.270 ;
        RECT 0.000 331.640 6.000 332.690 ;
        RECT 295.300 331.825 301.300 332.875 ;
        RECT 0.000 330.940 3.555 331.640 ;
        RECT 297.750 330.825 301.300 331.825 ;
        RECT 0.000 326.630 3.555 327.330 ;
        RECT 297.755 327.210 301.300 327.315 ;
        RECT 297.750 326.815 301.300 327.210 ;
        RECT 0.000 325.580 6.000 326.630 ;
        RECT 295.300 325.765 301.300 326.815 ;
        RECT 0.000 324.880 3.555 325.580 ;
        RECT 297.750 324.765 301.300 325.765 ;
        RECT 0.000 320.570 3.555 321.270 ;
        RECT 297.755 321.150 301.300 321.255 ;
        RECT 297.750 320.755 301.300 321.150 ;
        RECT 0.000 319.520 6.000 320.570 ;
        RECT 295.300 319.705 301.300 320.755 ;
        RECT 0.000 318.820 3.555 319.520 ;
        RECT 297.750 318.705 301.300 319.705 ;
        RECT 0.000 314.510 3.555 315.210 ;
        RECT 297.755 315.090 301.300 315.195 ;
        RECT 297.750 314.695 301.300 315.090 ;
        RECT 0.000 313.460 6.000 314.510 ;
        RECT 295.300 313.645 301.300 314.695 ;
        RECT 0.000 312.760 3.555 313.460 ;
        RECT 297.750 312.645 301.300 313.645 ;
        RECT 0.000 308.450 3.555 309.150 ;
        RECT 297.750 308.635 301.300 309.135 ;
        RECT 0.000 307.400 6.000 308.450 ;
        RECT 295.300 307.585 301.300 308.635 ;
        RECT 0.000 306.700 3.555 307.400 ;
        RECT 297.750 306.685 301.300 307.585 ;
        RECT 0.000 302.390 3.555 303.090 ;
        RECT 297.750 302.575 301.300 303.075 ;
        RECT 0.000 301.340 6.000 302.390 ;
        RECT 295.300 301.525 301.300 302.575 ;
        RECT 0.000 300.640 3.555 301.340 ;
        RECT 297.750 300.625 301.300 301.525 ;
        RECT 0.000 296.330 3.555 297.030 ;
        RECT 297.750 296.515 301.300 297.015 ;
        RECT 0.000 295.280 6.000 296.330 ;
        RECT 295.300 295.465 301.300 296.515 ;
        RECT 0.000 294.580 3.555 295.280 ;
        RECT 297.750 294.565 301.300 295.465 ;
        RECT 0.000 290.270 3.555 290.970 ;
        RECT 297.750 290.455 301.300 290.955 ;
        RECT 0.000 289.220 6.000 290.270 ;
        RECT 295.300 289.405 301.300 290.455 ;
        RECT 0.000 288.520 3.555 289.220 ;
        RECT 297.750 288.505 301.300 289.405 ;
        RECT 0.000 284.210 3.555 284.910 ;
        RECT 297.750 284.395 301.300 284.895 ;
        RECT 0.000 283.160 6.000 284.210 ;
        RECT 295.300 283.345 301.300 284.395 ;
        RECT 0.000 282.460 3.555 283.160 ;
        RECT 297.750 282.445 301.300 283.345 ;
        RECT 0.000 278.150 3.555 278.850 ;
        RECT 297.750 278.335 301.300 278.835 ;
        RECT 0.000 277.100 6.000 278.150 ;
        RECT 295.300 277.285 301.300 278.335 ;
        RECT 0.000 276.400 3.555 277.100 ;
        RECT 297.750 276.385 301.300 277.285 ;
        RECT 0.000 272.090 3.555 272.790 ;
        RECT 297.750 272.275 301.300 272.775 ;
        RECT 0.000 271.040 6.000 272.090 ;
        RECT 295.300 271.225 301.300 272.275 ;
        RECT 0.000 270.340 3.555 271.040 ;
        RECT 297.750 270.325 301.300 271.225 ;
        RECT 0.000 266.030 3.555 266.730 ;
        RECT 297.750 266.215 301.300 266.715 ;
        RECT 0.000 264.980 6.000 266.030 ;
        RECT 295.300 265.165 301.300 266.215 ;
        RECT 0.000 264.280 3.555 264.980 ;
        RECT 297.750 264.265 301.300 265.165 ;
        RECT 0.000 259.970 3.555 260.670 ;
        RECT 297.750 260.155 301.300 260.655 ;
        RECT 0.000 258.920 6.000 259.970 ;
        RECT 295.300 259.105 301.300 260.155 ;
        RECT 0.000 258.220 3.555 258.920 ;
        RECT 297.750 258.205 301.300 259.105 ;
        RECT 0.000 253.910 3.555 254.610 ;
        RECT 297.750 254.095 301.300 254.595 ;
        RECT 0.000 252.860 6.000 253.910 ;
        RECT 295.300 253.045 301.300 254.095 ;
        RECT 0.000 252.160 3.555 252.860 ;
        RECT 297.750 252.145 301.300 253.045 ;
        RECT 0.000 247.850 3.555 248.550 ;
        RECT 297.750 248.035 301.300 248.535 ;
        RECT 0.000 246.800 6.000 247.850 ;
        RECT 295.300 246.985 301.300 248.035 ;
        RECT 0.000 246.100 3.555 246.800 ;
        RECT 297.750 246.085 301.300 246.985 ;
        RECT 0.000 241.790 3.555 242.490 ;
        RECT 297.750 241.975 301.300 242.475 ;
        RECT 0.000 240.740 6.000 241.790 ;
        RECT 295.300 240.925 301.300 241.975 ;
        RECT 0.000 240.040 3.555 240.740 ;
        RECT 297.750 240.025 301.300 240.925 ;
        RECT 0.000 235.730 3.555 236.430 ;
        RECT 297.750 235.915 301.300 236.415 ;
        RECT 0.000 234.680 6.000 235.730 ;
        RECT 295.300 234.865 301.300 235.915 ;
        RECT 0.000 233.980 3.555 234.680 ;
        RECT 297.750 233.965 301.300 234.865 ;
        RECT 0.000 229.670 3.555 230.370 ;
        RECT 297.750 229.855 301.300 230.355 ;
        RECT 0.000 228.620 6.000 229.670 ;
        RECT 295.300 228.805 301.300 229.855 ;
        RECT 0.000 227.920 3.555 228.620 ;
        RECT 297.750 227.905 301.300 228.805 ;
        RECT 0.000 223.610 3.555 224.310 ;
        RECT 297.750 223.795 301.300 224.295 ;
        RECT 0.000 222.560 6.000 223.610 ;
        RECT 295.300 222.745 301.300 223.795 ;
        RECT 0.000 221.860 3.555 222.560 ;
        RECT 297.750 221.845 301.300 222.745 ;
        RECT 0.000 217.550 3.555 218.250 ;
        RECT 297.750 217.735 301.300 218.235 ;
        RECT 0.000 216.500 6.000 217.550 ;
        RECT 295.300 216.685 301.300 217.735 ;
        RECT 0.000 215.800 3.555 216.500 ;
        RECT 297.750 215.785 301.300 216.685 ;
        RECT 0.000 211.490 3.555 212.190 ;
        RECT 297.750 211.675 301.300 212.175 ;
        RECT 0.000 210.440 6.000 211.490 ;
        RECT 295.300 210.625 301.300 211.675 ;
        RECT 0.000 209.740 3.555 210.440 ;
        RECT 297.750 209.725 301.300 210.625 ;
        RECT 0.000 205.430 3.555 206.130 ;
        RECT 297.750 205.615 301.300 206.115 ;
        RECT 0.000 204.380 6.000 205.430 ;
        RECT 295.300 204.565 301.300 205.615 ;
        RECT 0.000 203.680 3.555 204.380 ;
        RECT 297.750 203.665 301.300 204.565 ;
        RECT 0.000 199.370 3.555 200.070 ;
        RECT 297.750 199.555 301.300 200.055 ;
        RECT 0.000 198.320 6.000 199.370 ;
        RECT 295.300 198.505 301.300 199.555 ;
        RECT 0.000 197.620 3.555 198.320 ;
        RECT 297.750 197.605 301.300 198.505 ;
        RECT 0.000 193.310 3.555 194.010 ;
        RECT 297.750 193.495 301.300 193.995 ;
        RECT 0.000 192.260 6.000 193.310 ;
        RECT 295.300 192.445 301.300 193.495 ;
        RECT 0.000 191.560 3.555 192.260 ;
        RECT 297.750 191.545 301.300 192.445 ;
        RECT 0.000 187.250 3.555 187.950 ;
        RECT 297.750 187.435 301.300 187.935 ;
        RECT 0.000 186.200 6.000 187.250 ;
        RECT 295.300 186.385 301.300 187.435 ;
        RECT 0.000 185.500 3.555 186.200 ;
        RECT 297.750 185.485 301.300 186.385 ;
        RECT 0.000 181.190 3.555 181.890 ;
        RECT 297.750 181.375 301.300 181.875 ;
        RECT 0.000 180.140 6.000 181.190 ;
        RECT 295.300 180.325 301.300 181.375 ;
        RECT 0.000 179.440 3.555 180.140 ;
        RECT 297.750 179.425 301.300 180.325 ;
        RECT 0.000 175.130 3.555 175.830 ;
        RECT 297.750 175.315 301.300 175.815 ;
        RECT 0.000 174.080 6.000 175.130 ;
        RECT 295.300 174.265 301.300 175.315 ;
        RECT 0.000 173.380 3.555 174.080 ;
        RECT 297.750 173.365 301.300 174.265 ;
        RECT 0.000 169.070 3.555 169.770 ;
        RECT 297.750 169.255 301.300 169.755 ;
        RECT 0.000 168.020 6.000 169.070 ;
        RECT 295.300 168.205 301.300 169.255 ;
        RECT 0.000 167.320 3.555 168.020 ;
        RECT 297.750 167.305 301.300 168.205 ;
        RECT 0.000 163.010 3.555 163.710 ;
        RECT 297.750 163.195 301.300 163.695 ;
        RECT 0.000 161.960 6.000 163.010 ;
        RECT 295.300 162.145 301.300 163.195 ;
        RECT 0.000 161.260 3.555 161.960 ;
        RECT 297.750 161.245 301.300 162.145 ;
        RECT 0.000 156.950 3.555 157.650 ;
        RECT 297.750 157.135 301.300 157.635 ;
        RECT 0.000 155.900 6.000 156.950 ;
        RECT 295.300 156.085 301.300 157.135 ;
        RECT 0.000 155.200 3.555 155.900 ;
        RECT 297.750 155.185 301.300 156.085 ;
        RECT 0.000 150.890 3.555 151.590 ;
        RECT 297.750 151.075 301.300 151.575 ;
        RECT 0.000 149.840 6.000 150.890 ;
        RECT 295.300 150.025 301.300 151.075 ;
        RECT 0.000 149.140 3.555 149.840 ;
        RECT 297.750 149.125 301.300 150.025 ;
        RECT 0.000 144.830 3.555 145.530 ;
        RECT 297.750 145.015 301.300 145.515 ;
        RECT 0.000 143.780 6.000 144.830 ;
        RECT 295.300 143.965 301.300 145.015 ;
        RECT 0.000 143.080 3.555 143.780 ;
        RECT 297.750 143.065 301.300 143.965 ;
        RECT 0.000 138.770 3.555 139.470 ;
        RECT 297.750 138.955 301.300 139.455 ;
        RECT 0.000 137.720 6.000 138.770 ;
        RECT 295.300 137.905 301.300 138.955 ;
        RECT 0.000 137.020 3.555 137.720 ;
        RECT 297.750 137.005 301.300 137.905 ;
        RECT 0.000 132.710 3.555 133.410 ;
        RECT 297.750 132.895 301.300 133.395 ;
        RECT 0.000 131.660 6.000 132.710 ;
        RECT 295.300 131.845 301.300 132.895 ;
        RECT 0.000 130.960 3.555 131.660 ;
        RECT 297.750 130.945 301.300 131.845 ;
        RECT 0.000 126.650 3.555 127.350 ;
        RECT 297.755 127.190 301.300 127.335 ;
        RECT 297.750 126.835 301.300 127.190 ;
        RECT 0.000 125.600 6.000 126.650 ;
        RECT 295.300 125.785 301.300 126.835 ;
        RECT 0.000 124.900 3.555 125.600 ;
        RECT 297.750 124.885 301.300 125.785 ;
        RECT 0.000 120.590 3.555 121.290 ;
        RECT 297.755 121.080 301.300 121.275 ;
        RECT 297.750 120.775 301.300 121.080 ;
        RECT 0.000 119.540 6.000 120.590 ;
        RECT 295.300 119.725 301.300 120.775 ;
        RECT 0.000 118.840 3.555 119.540 ;
        RECT 297.750 118.825 301.300 119.725 ;
        RECT 0.010 114.115 6.000 114.360 ;
        RECT 0.000 113.660 6.000 114.115 ;
        RECT 295.300 113.660 301.300 114.360 ;
        RECT 0.000 113.025 3.555 113.660 ;
        RECT 297.750 113.025 301.300 113.660 ;
        RECT 0.000 111.350 6.000 113.025 ;
        RECT 0.010 111.345 6.000 111.350 ;
        RECT 295.300 111.345 301.300 113.025 ;
        RECT 0.000 93.825 3.545 93.830 ;
        RECT 297.750 93.825 301.300 93.830 ;
        RECT 0.000 86.895 6.000 93.825 ;
        RECT 0.010 86.890 6.000 86.895 ;
        RECT 295.300 86.890 301.300 93.825 ;
        RECT 295.300 86.830 295.500 86.890 ;
        RECT 0.000 72.855 0.700 72.860 ;
        RECT 297.755 72.855 301.300 72.860 ;
        RECT 0.000 71.265 6.000 72.855 ;
        RECT 295.300 71.265 301.300 72.855 ;
        RECT 0.000 69.355 3.555 71.265 ;
        RECT 297.755 70.860 301.300 71.265 ;
        RECT 297.750 69.355 301.300 70.860 ;
        RECT 0.000 47.950 6.000 57.210 ;
        RECT 295.300 47.950 301.300 57.210 ;
        RECT 297.750 38.225 301.300 38.230 ;
        RECT 0.000 33.615 6.000 38.225 ;
        RECT 295.300 33.615 301.300 38.225 ;
        RECT 0.000 23.645 6.000 25.465 ;
        RECT 295.300 23.645 301.300 25.465 ;
        RECT 0.000 23.315 3.565 23.645 ;
        RECT 297.745 23.315 301.300 23.645 ;
        RECT 0.000 21.325 3.555 23.315 ;
        RECT 297.750 21.325 301.300 23.315 ;
        RECT 0.000 19.810 6.000 21.325 ;
        RECT 295.300 19.810 301.300 21.325 ;
        RECT 0.000 13.195 0.700 13.200 ;
        RECT 0.000 11.965 6.000 13.195 ;
        RECT 295.300 11.965 301.300 13.195 ;
        RECT 0.000 9.985 3.545 11.965 ;
        RECT 297.805 9.985 301.300 11.965 ;
        RECT 0.000 8.740 6.000 9.985 ;
        RECT 295.300 8.750 301.300 9.985 ;
        RECT 295.300 8.745 298.065 8.750 ;
        RECT 16.245 0.000 19.745 3.260 ;
        RECT 33.045 0.000 36.545 3.260 ;
        RECT 54.045 0.000 57.545 3.260 ;
        RECT 70.845 0.000 74.345 3.260 ;
        RECT 109.630 0.000 113.130 3.260 ;
        RECT 115.575 0.000 119.075 3.260 ;
        RECT 121.905 0.000 125.405 3.260 ;
        RECT 133.095 0.000 136.595 3.260 ;
        RECT 144.315 0.000 147.815 3.260 ;
        RECT 152.715 0.000 156.215 3.260 ;
        RECT 161.115 0.000 164.615 3.260 ;
        RECT 179.315 0.000 182.815 3.260 ;
        RECT 183.670 0.000 187.170 3.260 ;
        RECT 223.760 0.000 227.260 3.260 ;
        RECT 240.560 0.000 244.060 3.260 ;
        RECT 261.560 0.000 265.060 3.260 ;
        RECT 278.360 0.000 281.860 3.260 ;
    END
  END VSS
  PIN WEN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal1 ;
        RECT 288.510 5.985 289.140 5.990 ;
        RECT 288.510 5.955 289.420 5.985 ;
        RECT 288.510 5.695 290.025 5.955 ;
        RECT 288.510 5.685 289.420 5.695 ;
        RECT 288.510 5.650 289.140 5.685 ;
        RECT 288.655 5.200 288.995 5.265 ;
        RECT 288.430 4.800 289.220 5.200 ;
        RECT 288.655 4.735 288.995 4.800 ;
      LAYER Metal2 ;
        RECT 288.430 0.000 289.215 5.995 ;
    END
  END WEN[7]
  PIN WEN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal1 ;
        RECT 253.790 5.985 254.350 5.995 ;
        RECT 253.285 5.965 254.350 5.985 ;
        RECT 253.185 5.705 254.355 5.965 ;
        RECT 253.285 5.695 254.350 5.705 ;
        RECT 253.285 5.645 253.915 5.695 ;
        RECT 253.405 5.200 253.745 5.265 ;
        RECT 253.180 4.800 253.970 5.200 ;
        RECT 253.405 4.735 253.745 4.800 ;
      LAYER Metal2 ;
        RECT 253.205 0.000 253.985 6.000 ;
    END
  END WEN[6]
  PIN WEN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal1 ;
        RECT 249.780 5.950 250.340 5.980 ;
        RECT 250.710 5.950 251.340 5.985 ;
        RECT 249.775 5.690 251.340 5.950 ;
        RECT 249.780 5.680 250.340 5.690 ;
        RECT 250.710 5.645 251.340 5.690 ;
        RECT 250.855 5.200 251.195 5.265 ;
        RECT 250.630 4.800 251.420 5.200 ;
        RECT 250.855 4.735 251.195 4.800 ;
      LAYER Metal2 ;
        RECT 250.630 0.000 251.410 6.000 ;
    END
  END WEN[5]
  PIN WEN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal1 ;
        RECT 214.710 5.960 215.270 5.990 ;
        RECT 214.105 5.950 215.275 5.960 ;
        RECT 214.105 5.940 216.880 5.950 ;
        RECT 214.105 5.700 217.110 5.940 ;
        RECT 214.320 5.690 217.110 5.700 ;
        RECT 216.480 5.600 217.110 5.690 ;
        RECT 216.525 5.505 216.880 5.600 ;
        RECT 216.645 5.200 216.985 5.265 ;
        RECT 216.420 4.800 217.210 5.200 ;
        RECT 216.645 4.735 216.985 4.800 ;
      LAYER Metal2 ;
        RECT 216.400 0.000 217.185 5.955 ;
    END
  END WEN[4]
  PIN WEN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal1 ;
        RECT 81.990 5.975 82.620 5.990 ;
        RECT 83.305 5.975 83.865 5.980 ;
        RECT 81.950 5.950 84.110 5.975 ;
        RECT 81.950 5.690 84.470 5.950 ;
        RECT 81.950 5.670 84.110 5.690 ;
        RECT 81.990 5.650 82.620 5.670 ;
        RECT 82.100 5.260 82.440 5.325 ;
        RECT 81.875 4.860 82.665 5.260 ;
        RECT 82.100 4.795 82.440 4.860 ;
      LAYER Metal2 ;
        RECT 81.910 0.000 82.695 6.000 ;
    END
  END WEN[3]
  PIN WEN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal1 ;
        RECT 45.915 5.940 46.545 5.990 ;
        RECT 48.235 5.960 48.795 5.990 ;
        RECT 47.630 5.940 48.800 5.960 ;
        RECT 45.915 5.700 48.800 5.940 ;
        RECT 45.915 5.690 48.795 5.700 ;
        RECT 45.915 5.665 48.390 5.690 ;
        RECT 45.915 5.650 46.545 5.665 ;
        RECT 45.930 5.260 46.270 5.325 ;
        RECT 45.705 4.860 46.495 5.260 ;
        RECT 45.930 4.795 46.270 4.860 ;
      LAYER Metal2 ;
        RECT 45.685 5.650 46.545 5.990 ;
        RECT 45.685 0.000 46.470 5.650 ;
    END
  END WEN[2]
  PIN WEN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal1 ;
        RECT 44.190 5.980 44.820 5.990 ;
        RECT 44.190 5.950 45.035 5.980 ;
        RECT 44.190 5.690 45.640 5.950 ;
        RECT 44.190 5.680 45.035 5.690 ;
        RECT 44.190 5.665 44.945 5.680 ;
        RECT 44.190 5.650 44.820 5.665 ;
        RECT 44.385 5.260 44.725 5.325 ;
        RECT 44.160 4.860 44.950 5.260 ;
        RECT 44.385 4.795 44.725 4.860 ;
      LAYER Metal2 ;
        RECT 44.110 0.000 44.895 5.995 ;
    END
  END WEN[1]
  PIN WEN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    ANTENNADIFFAREA 0.490250 ;
    PORT
      LAYER Metal1 ;
        RECT 8.800 5.650 10.850 6.000 ;
        RECT 10.215 5.645 10.845 5.650 ;
        RECT 10.330 5.260 10.670 5.325 ;
        RECT 10.105 4.860 10.895 5.260 ;
        RECT 10.330 4.795 10.670 4.860 ;
      LAYER Metal2 ;
        RECT 10.215 5.980 10.845 5.985 ;
        RECT 10.085 0.000 10.870 5.980 ;
    END
  END WEN[0]
  PIN A[9]
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 99.650 0.000 100.435 6.000 ;
    END
  END A[9]
  OBS
      LAYER Nwell ;
        RECT 6.305 6.000 295.010 509.810 ;
      LAYER Metal1 ;
        RECT 6.000 6.000 295.300 509.810 ;
      LAYER Metal2 ;
        RECT 6.000 6.000 295.300 509.810 ;
      LAYER Metal3 ;
        RECT 6.000 83.900 295.300 509.810 ;
        RECT 6.000 83.145 295.500 83.900 ;
        RECT 6.000 82.675 295.300 83.145 ;
        RECT 6.000 81.920 295.500 82.675 ;
        RECT 6.000 6.000 295.300 81.920 ;
  END
END gf180mcu_ocd_ip_sram__sram1024x8m8wm1
END LIBRARY

