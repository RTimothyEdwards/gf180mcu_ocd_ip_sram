magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -1815 248 1815 275
rect -1815 -248 -1790 248
rect 1790 -248 1815 248
rect -1815 -275 1815 -248
<< via2 >>
rect -1790 -248 1790 248
<< metal3 >>
rect -1815 248 1815 275
rect -1815 -248 -1790 248
rect 1790 -248 1815 248
rect -1815 -275 1815 -248
<< end >>
