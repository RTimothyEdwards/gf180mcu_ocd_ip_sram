magic
tech gf180mcuD
magscale 1 10
timestamp 1763482574
<< error_s >>
rect 19225 65306 19230 65311
rect 19271 25190 19276 65306
rect 39909 25190 39915 65311
rect 19209 24246 19236 24302
rect 19225 24240 19230 24246
rect 19265 23908 19292 24246
<< psubdiff >>
rect 18967 25183 20040 65408
rect 39151 25183 40172 65718
rect 59602 745 59871 65715
<< metal1 >>
rect 0 623 700 65686
<< metal2 >>
rect 296 623 996 65693
<< metal3 >>
rect 296 341 996 1562
use M1_PSUB4310591302043_512x8m81  M1_PSUB4310591302043_512x8m81_0
timestamp 1763482574
transform -1 0 59970 0 1 65401
box 171 -29 59921 289
use M1_PSUB4310591302043_512x8m81  M1_PSUB4310591302043_512x8m81_1
timestamp 1763482574
transform -1 0 59970 0 1 775
box 171 -29 59921 289
use M1_PSUB4310591302044_512x8m81  M1_PSUB4310591302044_512x8m81_0
timestamp 1763476864
transform 1 0 59631 0 1 798
box -29 266 240 64574
use M1_PSUB4310591302044_512x8m81  M1_PSUB4310591302044_512x8m81_1
timestamp 1763476864
transform 1 0 18997 0 1 798
box -29 266 240 64574
use M1_PSUB4310591302044_512x8m81  M1_PSUB4310591302044_512x8m81_2
timestamp 1763476864
transform 1 0 39932 0 1 798
box -29 266 240 64574
use M1_PSUB4310591302044_512x8m81  M1_PSUB4310591302044_512x8m81_3
timestamp 1763476864
transform 1 0 78 0 1 798
box -29 266 240 64574
use M1_PSUB4310591302045_512x8m81  M1_PSUB4310591302045_512x8m81_0
timestamp 1763476864
transform 1 0 39286 0 1 25213
box -29 -29 589 40099
use M1_PSUB4310591302045_512x8m81  M1_PSUB4310591302045_512x8m81_1
timestamp 1763476864
transform 1 0 19294 0 1 25213
box -29 -29 589 40099
use M1_PSUB4310591302046_512x8m81  M1_PSUB4310591302046_512x8m81_0
timestamp 1763476864
transform 1 0 19294 0 1 23937
box -29 -29 20539 309
<< labels >>
flabel metal3 s 646 465 646 465 0 FreeSans 313 0 0 0 VDD
port 1 nsew
<< properties >>
string path 4.620 11.160 4.620 0.000 
<< end >>
