magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< psubdiff >>
rect -996 23 996 57
rect -996 -23 -963 23
rect 963 -23 996 23
rect -996 -58 996 -23
<< psubdiffcont >>
rect -963 -23 963 23
<< metal1 >>
rect -990 23 990 51
rect -990 -23 -963 23
rect 963 -23 990 23
rect -990 -51 990 -23
<< end >>
