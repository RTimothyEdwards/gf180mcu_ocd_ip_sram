magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< psubdiff >>
rect -2018 787 2018 800
rect -2018 -787 -2005 787
rect 2005 -787 2018 787
rect -2018 -800 2018 -787
<< psubdiffcont >>
rect -2005 -787 2005 787
<< metal1 >>
rect -2013 787 2013 795
rect -2013 -787 -2005 787
rect 2005 -787 2013 787
rect -2013 -795 2013 -787
<< end >>
