magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -487 257 487 275
rect -487 -257 -471 257
rect 471 -257 487 257
rect -487 -275 487 -257
<< via2 >>
rect -471 -257 471 257
<< metal3 >>
rect -487 257 487 275
rect -487 -257 -471 257
rect 471 -257 487 257
rect -487 -275 487 -257
<< end >>
