magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< nwell >>
rect -328 -58 14 320
rect 15 -58 337 320
rect -328 -66 337 -58
rect 338 -66 667 320
rect 668 -66 986 320
rect 987 -66 1342 320
<< polysilicon >>
rect -266 253 -211 288
rect -106 253 -50 288
rect 55 253 111 288
rect 215 253 271 288
rect 376 253 432 288
rect 536 253 592 288
rect 697 253 753 288
rect 857 253 913 288
rect 1018 253 1074 288
rect 1178 253 1234 288
rect -266 -34 -211 0
rect -106 -34 -50 0
rect 55 -34 111 0
rect 215 -34 271 0
rect 376 -34 432 0
rect 536 -34 592 0
rect 697 -34 753 0
rect 857 -34 913 0
rect 1018 -34 1074 0
rect 1178 -34 1234 0
use pmos_5p04310591302030_512x8m81  pmos_5p04310591302030_512x8m81_0
timestamp 1763564386
transform 1 0 -14 0 1 0
box -426 -86 1422 339
<< end >>
