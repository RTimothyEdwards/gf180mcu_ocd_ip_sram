magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal1 >>
rect -45 18 487 46
rect -45 -170 -18 18
rect 461 -170 487 18
rect -45 -198 487 -170
<< via1 >>
rect -18 -170 461 18
<< metal2 >>
rect -45 18 487 46
rect -45 -170 -18 18
rect 461 -170 487 18
rect -45 -198 487 -170
<< end >>
