magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< error_s >>
rect 0 74 65 88
rect 0 17 3 74
rect 0 0 65 17
use via1_R90_3v1024x8m81_0  via1_R90_3v1024x8m81_0_0
timestamp 1764525316
transform 1 0 0 0 1 0
box 0 0 65 89
use via2_R90_3v1024x8m81_0  via2_R90_3v1024x8m81_0_0
timestamp 1764525316
transform 1 0 0 0 1 0
box 0 0 65 89
<< end >>
