magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< nwell >>
rect -174 -86 230 1504
<< pmos >>
rect 0 0 56 1418
<< pdiff >>
rect -88 1405 0 1418
rect -88 13 -75 1405
rect -29 13 0 1405
rect -88 0 0 13
rect 56 1405 144 1418
rect 56 13 85 1405
rect 131 13 144 1405
rect 56 0 144 13
<< pdiffc >>
rect -75 13 -29 1405
rect 85 13 131 1405
<< polysilicon >>
rect 0 1418 56 1462
rect 0 -44 56 0
<< metal1 >>
rect -75 1405 -29 1418
rect -75 0 -29 13
rect 85 1405 131 1418
rect 85 0 131 13
<< labels >>
flabel pdiffc -40 709 -40 709 0 FreeSans 186 0 0 0 S
flabel pdiffc 96 709 96 709 0 FreeSans 186 0 0 0 D
<< end >>
