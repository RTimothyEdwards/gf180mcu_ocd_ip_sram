magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< nwell >>
rect -202 -86 362 404
<< pmos >>
rect -28 0 28 318
rect 132 0 188 318
<< pdiff >>
rect -116 281 -28 318
rect -116 13 -103 281
rect -57 13 -28 281
rect -116 0 -28 13
rect 28 281 132 318
rect 28 13 57 281
rect 103 13 132 281
rect 28 0 132 13
rect 188 281 276 318
rect 188 13 217 281
rect 263 13 276 281
rect 188 0 276 13
<< pdiffc >>
rect -103 13 -57 281
rect 57 13 103 281
rect 217 13 263 281
<< polysilicon >>
rect -28 318 28 362
rect 132 318 188 362
rect -28 -44 28 0
rect 132 -44 188 0
<< metal1 >>
rect -103 281 -57 318
rect -103 0 -57 13
rect 57 281 103 318
rect 57 0 103 13
rect 217 281 263 318
rect 217 0 263 13
<< labels >>
flabel pdiffc 80 159 80 159 0 FreeSans 186 0 0 0 D
flabel pdiffc -68 159 -68 159 0 FreeSans 186 0 0 0 S
flabel pdiffc 228 159 228 159 0 FreeSans 186 0 0 0 S
<< end >>
