magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nwell >>
rect 3206 1787 3623 1813
rect 2608 1701 3623 1787
rect 1508 1611 3623 1701
rect -372 851 3623 1611
rect -372 837 3206 851
rect 3456 850 3493 851
rect -123 795 3206 837
rect -123 767 1078 795
<< pdiff >>
rect 1969 1491 2053 1603
<< polysilicon >>
rect 2826 1866 3286 1918
rect 1849 1695 1905 1800
rect 2141 1711 2197 1778
rect 2599 1775 2966 1817
rect 1697 1652 1946 1695
rect 2141 1652 2395 1711
rect 1697 1643 1753 1652
rect 1857 1643 1913 1652
rect 2141 1645 2197 1652
rect 2750 1505 2806 1775
rect 2910 1505 2966 1775
rect 3070 1504 3126 1866
rect 3230 1504 3286 1866
rect 1750 1256 2207 1313
rect 1750 1255 1967 1256
rect 1750 1146 1806 1255
rect 1911 1146 1967 1255
rect 2071 1255 2207 1256
rect 2071 1248 2151 1255
rect 2071 1146 2127 1248
rect 2384 1237 2440 1417
rect 64 816 120 832
rect 224 816 280 832
rect 386 816 442 832
rect 546 816 602 832
rect 707 816 763 832
rect 867 816 923 832
rect 64 757 1050 816
rect 64 711 120 757
rect 224 711 280 757
rect 385 711 441 757
rect 545 711 601 757
rect 706 711 762 757
rect 866 711 922 757
rect 1155 561 1211 855
rect 1444 793 1500 858
rect 1418 721 1500 793
rect 1444 570 1500 721
rect 2384 695 2440 943
rect 2752 808 3004 815
rect 2752 762 3114 808
rect 2752 743 2968 762
rect 2752 713 2808 743
rect 2912 698 2968 743
rect 1155 276 1211 343
rect 1444 331 1500 344
rect 1750 296 2326 338
rect 2384 296 2440 524
rect 3072 188 3128 365
rect 3232 188 3288 365
rect 3072 116 3288 188
<< metal1 >>
rect 1948 1997 2058 2214
rect 1948 1944 2463 1997
rect 135 1165 217 1404
rect 449 1165 530 1404
rect 772 1195 819 1404
rect 1517 1198 1563 1899
rect 1780 1346 1827 1929
rect 1948 1799 2100 1944
rect 2201 1733 2282 1889
rect 2412 1822 2463 1944
rect 1880 1681 2282 1733
rect 1982 1402 2061 1617
rect 2201 1506 2282 1681
rect 2339 1603 2516 1711
rect 2675 1666 3362 1715
rect 2675 1462 2721 1666
rect 2995 1452 3041 1666
rect 3315 1584 3362 1666
rect 3315 1452 3361 1584
rect 2168 1350 2521 1402
rect 1667 1262 2062 1346
rect 786 1165 819 1195
rect -11 816 35 1012
rect 311 816 357 1012
rect 630 816 677 1011
rect 943 816 993 1012
rect -11 732 993 816
rect -11 545 35 732
rect 135 243 217 630
rect 311 545 357 732
rect 449 243 530 630
rect 630 545 677 732
rect 763 243 844 630
rect 943 545 993 732
rect 1240 787 1286 920
rect 1240 727 1336 787
rect 1240 521 1286 727
rect 1528 476 1575 922
rect 1667 380 1748 1262
rect 1824 330 1905 1205
rect 1981 380 2062 1262
rect 2168 1260 2219 1350
rect 2137 330 2219 1206
rect 2298 604 2352 1262
rect 2837 669 2883 996
rect 1512 180 1559 327
rect 1824 247 2219 330
rect 2297 564 2352 604
rect 2297 302 2347 564
rect 2694 273 2745 484
rect 2997 273 3044 444
rect 3311 273 3363 452
rect 2694 227 3363 273
rect 1512 178 2629 180
rect 1512 133 3183 178
rect 2571 132 3183 133
<< metal2 >>
rect 2153 1638 2410 1706
rect 1982 1402 2061 1617
rect 2153 772 2219 1638
rect 2335 372 2398 1438
rect 2595 742 2661 1925
rect 3026 770 3092 1925
rect 2335 280 2402 372
<< metal3 >>
rect 1479 1858 3007 1923
rect -249 1051 3504 1618
rect 1043 774 2891 842
rect -249 -251 3519 669
use M1_NACTIVE4310591302038_256x8m81  M1_NACTIVE4310591302038_256x8m81_0
timestamp 1763766357
transform 1 0 3468 0 1 1365
box -36 -292 36 292
use M1_NACTIVE4310591302041_256x8m81  M1_NACTIVE4310591302041_256x8m81_0
timestamp 1763766357
transform 1 0 334 0 1 1373
box -490 -36 490 36
use M1_NWELL_01_R270_256x8m81  M1_NWELL_01_R270_256x8m81_0
timestamp 1763766357
transform 0 1 -217 -1 0 1110
box -273 -154 273 154
use M1_PACTIVE4310591302034_256x8m81  M1_PACTIVE4310591302034_256x8m81_0
timestamp 1763766357
transform 1 0 -217 0 1 508
box -36 -128 36 128
use M1_PACTIVE4310591302039_256x8m81  M1_PACTIVE4310591302039_256x8m81_0
timestamp 1763766357
transform 1 0 3468 0 1 -126
box -36 -95 36 95
use M1_PACTIVE4310591302040_256x8m81  M1_PACTIVE4310591302040_256x8m81_0
timestamp 1763766357
transform 1 0 478 0 1 236
box -522 -36 522 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_0
timestamp 1763766357
transform 0 -1 1070 1 0 780
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_1
timestamp 1763766357
transform 1 0 2475 0 1 328
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_2
timestamp 1763766357
transform 1 0 1910 0 1 1709
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_3
timestamp 1763766357
transform 1 0 2368 0 1 1682
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_4
timestamp 1763766357
transform 1 0 2178 0 1 1284
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_5
timestamp 1763766357
transform 1 0 2426 0 1 1382
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_6
timestamp 1763766357
transform 1 0 2629 0 1 1809
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_7
timestamp 1763766357
transform 1 0 2297 0 1 325
box -36 -36 36 36
use M1_POLY24310591302033_256x8m81  M1_POLY24310591302033_256x8m81_0
timestamp 1763766357
transform -1 0 1487 0 -1 298
box -62 -36 62 36
use M1_POLY24310591302033_256x8m81  M1_POLY24310591302033_256x8m81_1
timestamp 1763766357
transform -1 0 1359 0 -1 757
box -62 -36 62 36
use M1_POLY24310591302033_256x8m81  M1_POLY24310591302033_256x8m81_2
timestamp 1763766357
transform 1 0 2883 0 -1 1902
box -62 -36 62 36
use M1_POLY24310591302033_256x8m81  M1_POLY24310591302033_256x8m81_3
timestamp 1763766357
transform 1 0 3216 0 1 151
box -62 -36 62 36
use M1_POLY24310591302033_256x8m81  M1_POLY24310591302033_256x8m81_4
timestamp 1763766357
transform 1 0 1180 0 1 245
box -62 -36 62 36
use M1_POLY24310591302033_256x8m81  M1_POLY24310591302033_256x8m81_5
timestamp 1763766357
transform -1 0 3055 0 1 799
box -62 -36 62 36
use M1_PSUB_02_256x8m81  M1_PSUB_02_256x8m81_0
timestamp 1763766357
transform 1 0 2462 0 1 1873
box -56 -57 56 58
use M2_M1$$168351788_R90_256x8m81  M2_M1$$168351788_R90_256x8m81_0
timestamp 1763766357
transform 0 -1 2520 1 0 326
box -46 -119 46 118
use M2_M1$$168351788_R90_256x8m81  M2_M1$$168351788_R90_256x8m81_1
timestamp 1763766357
transform 0 -1 2402 1 0 1397
box -46 -119 46 118
use M2_M1431059130200_256x8m81  M2_M1431059130200_256x8m81_0
timestamp 1763766357
transform 1 0 1183 0 1 245
box -63 -34 63 34
use M2_M1431059130200_256x8m81  M2_M1431059130200_256x8m81_1
timestamp 1763766357
transform 1 0 1110 0 1 783
box -63 -34 63 34
use M2_M1431059130200_256x8m81  M2_M1431059130200_256x8m81_2
timestamp 1763766357
transform 1 0 2828 0 1 809
box -63 -34 63 34
use M2_M1431059130200_256x8m81  M2_M1431059130200_256x8m81_3
timestamp 1763766357
transform -1 0 3057 0 1 799
box -63 -34 63 34
use M3_M2431059130207_256x8m81  M3_M2431059130207_256x8m81_0
timestamp 1763766357
transform 1 0 2828 0 1 809
box -63 -35 63 35
use M3_M2431059130207_256x8m81  M3_M2431059130207_256x8m81_1
timestamp 1763766357
transform 1 0 1106 0 1 782
box -63 -35 63 35
use nmos_5p0431059130208_256x8m81  nmos_5p0431059130208_256x8m81_0
timestamp 1763766357
transform -1 0 2440 0 1 564
box -88 -44 144 133
use nmos_5p0431059130208_256x8m81  nmos_5p0431059130208_256x8m81_1
timestamp 1763766357
transform 1 0 1849 0 -1 1932
box -88 -44 144 133
use nmos_5p04310591302033_256x8m81  nmos_5p04310591302033_256x8m81_0
timestamp 1763766357
transform 1 0 2141 0 -1 1871
box -92 -44 148 100
use nmos_5p04310591302044_256x8m81  nmos_5p04310591302044_256x8m81_0
timestamp 1763766357
transform -1 0 1500 0 1 378
box -88 -44 144 249
use nmos_5p04310591302045_256x8m81  nmos_5p04310591302045_256x8m81_0
timestamp 1763766357
transform 1 0 3100 0 -1 669
box -116 -44 276 309
use nmos_5p04310591302045_256x8m81  nmos_5p04310591302045_256x8m81_1
timestamp 1763766357
transform 1 0 2780 0 -1 669
box -116 -44 276 309
use nmos_5p04310591302046_256x8m81  nmos_5p04310591302046_256x8m81_0
timestamp 1763766357
transform -1 0 782 0 -1 669
box -228 -44 806 241
use nmos_5p04310591302050_256x8m81  nmos_5p04310591302050_256x8m81_0
timestamp 1763766357
transform -1 0 2071 0 1 380
box -144 -44 409 255
use nmos_5p04310591302052_256x8m81  nmos_5p04310591302052_256x8m81_0
timestamp 1763766357
transform -1 0 1211 0 1 380
box -88 -44 144 193
use pmos_1p2$$171625516_256x8m81  pmos_1p2$$171625516_256x8m81_0
timestamp 1763766357
transform 1 0 1739 0 -1 1603
box -216 -86 348 192
use pmos_5p04310591302013_256x8m81  pmos_5p04310591302013_256x8m81_0
timestamp 1763766357
transform -1 0 2071 0 1 895
box -230 -86 495 297
use pmos_5p04310591302014_256x8m81  pmos_5p04310591302014_256x8m81_0
timestamp 1763766357
transform -1 0 2440 0 1 984
box -174 -86 230 297
use pmos_5p04310591302038_256x8m81  pmos_5p04310591302038_256x8m81_0
timestamp 1763766357
transform 1 0 2141 0 -1 1603
box -174 -86 230 198
use pmos_5p04310591302047_256x8m81  pmos_5p04310591302047_256x8m81_0
timestamp 1763766357
transform -1 0 1211 0 1 895
box -174 -86 230 459
use pmos_5p04310591302048_256x8m81  pmos_5p04310591302048_256x8m81_0
timestamp 1763766357
transform -1 0 1500 0 1 864
box -174 -86 230 506
use pmos_5p04310591302049_256x8m81  pmos_5p04310591302049_256x8m81_0
timestamp 1763766357
transform -1 0 783 0 1 866
box -314 -86 894 438
use pmos_5p04310591302051_256x8m81  pmos_5p04310591302051_256x8m81_0
timestamp 1763766357
transform 1 0 2778 0 1 935
box -202 -86 362 615
use pmos_5p04310591302051_256x8m81  pmos_5p04310591302051_256x8m81_1
timestamp 1763766357
transform 1 0 3098 0 1 935
box -202 -86 362 615
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_0
timestamp 1763766357
transform -1 0 2218 0 1 760
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_1
timestamp 1763766357
transform -1 0 1897 0 1 760
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_2
timestamp 1763766357
transform 0 -1 2958 1 0 1848
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_3
timestamp 1763766357
transform 0 -1 1724 1 0 1848
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_4
timestamp 1763766357
transform 1 0 3436 0 1 -238
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_5
timestamp 1763766357
transform 1 0 144 0 1 1052
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_6
timestamp 1763766357
transform 1 0 456 0 1 1052
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_7
timestamp 1763766357
transform 1 0 770 0 1 1052
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_8
timestamp 1763766357
transform 1 0 456 0 1 441
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_9
timestamp 1763766357
transform 1 0 144 0 1 441
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_10
timestamp 1763766357
transform 1 0 3157 0 1 1052
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_11
timestamp 1763766357
transform 1 0 3157 0 1 1402
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_12
timestamp 1763766357
transform 1 0 3158 0 1 441
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_13
timestamp 1763766357
transform 1 0 2467 0 1 1052
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_14
timestamp 1763766357
transform 1 0 2482 0 1 441
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_15
timestamp 1763766357
transform 1 0 771 0 1 441
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_16
timestamp 1763766357
transform 1 0 1912 0 1 1402
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_17
timestamp 1763766357
transform 1 0 1618 0 1 1402
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_18
timestamp 1763766357
transform 1 0 -249 0 1 1052
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_19
timestamp 1763766357
transform 1 0 -249 0 1 441
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_20
timestamp 1763766357
transform 1 0 3436 0 1 1052
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_21
timestamp 1763766357
transform 1 0 3436 0 1 1402
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_22
timestamp 1763766357
transform 1 0 1071 0 1 1052
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_23
timestamp 1763766357
transform 1 0 1346 0 1 1052
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_24
timestamp 1763766357
transform 1 0 1071 0 1 375
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_25
timestamp 1763766357
transform 1 0 1346 0 1 375
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_26
timestamp 1763766357
transform 1 0 2023 0 1 1402
box -9 0 73 215
use via1_R270_256x8m81  via1_R270_256x8m81_0
timestamp 1763766357
transform 0 1 2339 -1 0 1705
box 0 0 67 89
use via1_x2_256x8m81  via1_x2_256x8m81_0
timestamp 1763766357
transform -1 0 2660 0 1 1763
box -8 0 72 222
<< labels >>
rlabel metal3 s -149 450 -149 450 4 vss
port 1 nsew
rlabel metal3 s -178 1491 -178 1491 4 vdd
port 2 nsew
rlabel metal2 s 2633 1885 2633 1885 4 qp
port 3 nsew
rlabel metal2 s 3080 1885 3080 1885 4 qn
port 4 nsew
rlabel metal1 s 2539 328 2539 328 4 se
port 5 nsew
rlabel metal1 s 2457 1882 2457 1882 4 vss
port 1 nsew
rlabel metal1 s 1129 252 1129 252 4 GWE
port 7 nsew
rlabel metal1 s 321 801 321 801 4 q
port 6 nsew
<< properties >>
string path 21.660 12.815 21.660 12.970 
<< end >>
