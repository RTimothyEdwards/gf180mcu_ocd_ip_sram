magic
tech gf180mcuD
magscale 1 10
timestamp 1763485967
<< nwell >>
rect -41 8409 610 11860
rect -13 4474 627 4880
rect -130 4462 627 4474
rect -130 4019 609 4462
<< pmos >>
rect 172 10921 228 11239
rect 332 10921 388 11239
rect 172 10416 228 10733
rect 332 10416 388 10733
rect 67 4108 123 4247
rect 319 4108 375 4247
<< pdiff >>
rect 46 11195 172 11239
rect 46 11149 97 11195
rect 143 11149 172 11195
rect 46 11013 172 11149
rect 46 10967 97 11013
rect 143 10967 172 11013
rect 46 10921 172 10967
rect 228 11195 332 11239
rect 228 11149 257 11195
rect 303 11149 332 11195
rect 228 11013 332 11149
rect 228 10967 257 11013
rect 303 10967 332 11013
rect 228 10921 332 10967
rect 388 11195 523 11239
rect 388 11149 443 11195
rect 489 11149 523 11195
rect 388 11013 523 11149
rect 388 10967 443 11013
rect 489 10967 523 11013
rect 388 10921 523 10967
rect 46 10690 172 10733
rect 46 10644 97 10690
rect 143 10644 172 10690
rect 46 10508 172 10644
rect 46 10462 97 10508
rect 143 10462 172 10508
rect 46 10416 172 10462
rect 228 10690 332 10733
rect 228 10644 257 10690
rect 303 10644 332 10690
rect 228 10508 332 10644
rect 228 10462 257 10508
rect 303 10462 332 10508
rect 228 10416 332 10462
rect 388 10690 523 10733
rect 388 10644 443 10690
rect 489 10644 523 10690
rect 388 10508 523 10644
rect 388 10462 443 10508
rect 489 10462 523 10508
rect 388 10416 523 10462
rect -44 4202 67 4247
rect -44 4155 -24 4202
rect 22 4155 67 4202
rect -44 4108 67 4155
rect 123 4201 319 4247
rect 123 4155 208 4201
rect 254 4155 319 4201
rect 123 4108 319 4155
rect 375 4201 523 4247
rect 375 4155 447 4201
rect 493 4155 523 4201
rect 375 4108 523 4155
<< pdiffc >>
rect 97 11149 143 11195
rect 97 10967 143 11013
rect 257 11149 303 11195
rect 257 10967 303 11013
rect 443 11149 489 11195
rect 443 10967 489 11013
rect 97 10644 143 10690
rect 97 10462 143 10508
rect 257 10644 303 10690
rect 257 10462 303 10508
rect 443 10644 489 10690
rect 443 10462 489 10508
rect -24 4155 22 4202
rect 208 4155 254 4201
rect 447 4155 493 4201
<< nsubdiff >>
rect 119 11552 523 11712
<< polysilicon >>
rect 172 11239 228 11436
rect 332 11239 388 11436
rect 172 10733 228 10921
rect 332 10733 388 10921
rect 172 10352 228 10416
rect 332 10352 388 10416
rect 172 10268 388 10352
rect 218 10267 304 10268
rect 248 10119 304 10267
rect 250 8475 306 8555
rect 250 6866 306 7513
rect 250 5995 306 6152
rect 250 5641 306 5852
rect 67 4386 375 4485
rect 67 4247 123 4386
rect 319 4247 375 4386
rect 67 4083 123 4108
rect 67 4010 194 4083
rect 319 4072 375 4108
rect 138 3948 194 4010
rect 306 4010 375 4072
rect 306 3948 362 4010
rect 138 3781 194 3810
rect 306 3781 362 3810
<< metal1 >>
rect 49 11562 523 11717
rect 74 11434 494 11562
rect 74 11195 159 11434
rect 74 11149 97 11195
rect 143 11149 159 11195
rect 74 11013 159 11149
rect 74 10967 97 11013
rect 143 10967 159 11013
rect 74 10690 159 10967
rect 222 11195 337 11382
rect 222 11149 257 11195
rect 303 11149 337 11195
rect 222 11013 337 11149
rect 222 10967 257 11013
rect 303 10967 337 11013
rect 222 10930 337 10967
rect 402 11195 494 11434
rect 402 11149 443 11195
rect 489 11149 494 11195
rect 402 11013 494 11149
rect 402 10967 443 11013
rect 489 10967 494 11013
rect 74 10644 97 10690
rect 143 10644 159 10690
rect 74 10508 159 10644
rect 74 10462 97 10508
rect 143 10462 159 10508
rect 74 10425 159 10462
rect 222 10690 337 10879
rect 222 10644 257 10690
rect 303 10644 337 10690
rect 222 10508 337 10644
rect 222 10462 257 10508
rect 303 10462 337 10508
rect 222 10425 337 10462
rect 402 10690 494 10967
rect 402 10644 443 10690
rect 489 10644 494 10690
rect 402 10508 494 10644
rect 402 10462 443 10508
rect 489 10462 494 10508
rect 402 10425 494 10462
rect 68 9710 219 9890
rect 333 9710 494 9890
rect 119 9065 182 9231
rect 130 8751 182 9065
rect 119 8647 182 8751
rect 119 7557 189 8647
rect 236 8296 332 8479
rect 381 7478 445 9227
rect 45 7381 445 7478
rect 43 7103 523 7237
rect 113 6958 495 7055
rect 113 6191 188 6958
rect 380 6232 457 6816
rect 113 4967 181 6191
rect 239 5939 331 6074
rect 239 5773 331 5884
rect 378 4810 457 6232
rect -41 4675 31 4693
rect -41 4591 73 4675
rect -41 4202 31 4591
rect 198 4396 374 4493
rect -41 4155 -24 4202
rect 22 4155 31 4202
rect -41 4117 31 4155
rect 205 4201 288 4317
rect 205 4155 208 4201
rect 254 4155 288 4201
rect 37 3742 120 3971
rect 205 3851 288 4155
rect 443 4201 523 4693
rect 443 4155 447 4201
rect 493 4155 523 4201
rect 443 4117 523 4155
rect 378 3742 457 3971
rect 37 3470 457 3742
<< metal2 >>
rect 68 11314 124 11715
rect 216 11435 344 11717
rect 245 11434 344 11435
rect 68 11258 327 11314
rect 68 9109 124 11258
rect 438 10808 494 11715
rect 285 10752 494 10808
rect 248 7338 304 8406
rect 191 7282 304 7338
rect 191 6246 247 7282
rect 438 6957 494 10752
rect 143 6190 247 6246
rect 143 5838 199 6190
rect 411 6074 474 6873
rect 260 5977 474 6074
rect 143 5782 312 5838
rect 143 4317 199 5782
rect 411 5094 474 5977
rect 270 4997 474 5094
rect 270 4396 330 4997
rect 143 4137 290 4317
rect 172 3520 272 3749
<< metal3 >>
rect -65 10338 525 11716
rect -41 7007 525 8407
rect -41 6761 525 6901
rect -41 6519 525 6659
rect -41 6278 525 6418
rect -41 6036 525 6176
rect -41 5504 525 5644
rect -41 5262 525 5402
rect -41 5020 525 5160
rect -41 4778 525 4918
rect -41 4190 525 4632
rect -41 3519 525 3974
use M1_NWELL05_512x8m81  M1_NWELL05_512x8m81_0
timestamp 1763476864
transform 1 0 285 0 1 11632
box -265 -159 265 159
use M1_NWELL09_512x8m81  M1_NWELL09_512x8m81_1
timestamp 1763476864
transform 1 0 279 0 1 4633
box -320 -159 320 159
use M1_POLY24310591302030_512x8m81  M1_POLY24310591302030_512x8m81_0
timestamp 1763476864
transform 1 0 272 0 1 10310
box -95 -36 95 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1763476864
transform 1 0 253 0 1 4443
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1763476864
transform 1 0 290 0 1 5810
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_2
timestamp 1763476864
transform 1 0 281 0 1 6037
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_6
timestamp 1763476864
transform 1 0 276 0 1 8442
box -36 -36 36 36
use M1_PSUB$$45111340_512x8m81  M1_PSUB$$45111340_512x8m81_0
timestamp 1763476864
transform 1 0 120 0 1 7168
box -56 -58 56 58
use M1_PSUB$$45111340_512x8m81  M1_PSUB$$45111340_512x8m81_1
timestamp 1763476864
transform 1 0 435 0 1 7168
box -56 -58 56 58
use M1_PSUB$$47122476_512x8m81  M1_PSUB$$47122476_512x8m81_0
timestamp 1763476864
transform 1 0 269 0 1 3544
box -223 -58 254 57
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_0
timestamp 1763476864
transform 1 0 247 0 1 4227
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_2
timestamp 1763476864
transform 1 0 106 0 1 9800
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_3
timestamp 1763476864
transform 1 0 108 0 1 9168
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_4
timestamp 1763476864
transform 1 0 281 0 1 11285
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_5
timestamp 1763476864
transform 1 0 276 0 1 8389
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_6
timestamp 1763476864
transform 1 0 456 0 1 9800
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_7
timestamp 1763476864
transform 1 0 281 0 1 10780
box -34 -63 34 63
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_0
timestamp 1763476864
transform 1 0 304 0 1 4442
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_1
timestamp 1763476864
transform 1 0 295 0 1 5810
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_5
timestamp 1763476864
transform 0 1 117 -1 0 7429
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_6
timestamp 1763476864
transform 1 0 344 0 1 7162
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_9
timestamp 1763476864
transform 1 0 459 0 1 7004
box -35 -56 35 55
use M3_M2431059130201_512x8m81  M3_M2431059130201_512x8m81_1
timestamp 1763476864
transform 1 0 344 0 1 7157
box -35 -63 35 63
use nmos_1p2$$47119404_512x8m81  nmos_1p2$$47119404_512x8m81_1
timestamp 1763476864
transform 1 0 264 0 -1 6826
box -102 -44 130 679
use nmos_1p2$$47119404_512x8m81  nmos_1p2$$47119404_512x8m81_3
timestamp 1763476864
transform 1 0 264 0 -1 8190
box -102 -44 130 679
use nmos_5p0431059130202_512x8m81  nmos_5p0431059130202_512x8m81_0
timestamp 1763476864
transform 1 0 170 0 1 3853
box -124 -44 285 98
use pmos_1p2$$46889004_512x8m81  pmos_1p2$$46889004_512x8m81_1
timestamp 1763476864
transform 1 0 264 0 -1 5601
box -188 -86 216 721
use pmos_5p0431059130201_512x8m81  pmos_5p0431059130201_512x8m81_0
timestamp 1763476864
transform 1 0 248 0 -1 10077
box -174 -86 230 721
use pmos_5p0431059130201_512x8m81  pmos_5p0431059130201_512x8m81_1
timestamp 1763476864
transform 1 0 250 0 -1 9231
box -174 -86 230 721
use via1_2_512x8m81  via1_2_512x8m81_0
timestamp 1763476864
transform 1 0 174 0 1 3559
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_0
timestamp 1763476864
transform 1 0 259 0 1 5979
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_2
timestamp 1763476864
transform 0 -1 343 1 0 11435
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_3
timestamp 1763476864
transform 0 -1 343 1 0 11621
box 0 0 65 89
use via2_R90_512x8m81  via2_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 373 1 0 11435
box 0 0 65 89
use via2_R90_512x8m81  via2_R90_512x8m81_1
timestamp 1763476864
transform 0 -1 373 1 0 11621
box 0 0 65 89
<< labels >>
rlabel metal1 s 318 4597 318 4597 4 vdd
port 2 nsew
rlabel metal1 s 229 10312 229 10312 4 pcb
port 8 nsew
rlabel metal2 s 105 11421 105 11421 4 bb
port 4 nsew
rlabel metal2 s 428 11421 428 11421 4 b
port 3 nsew
rlabel metal3 s 303 6306 303 6306 4 vss
port 1 nsew
rlabel metal3 s 318 11384 318 11384 4 vdd
port 2 nsew
rlabel metal2 s 281 4463 281 4463 4 ypass
port 6 nsew
rlabel metal1 s 450 5046 450 5046 4 d
port 7 nsew
<< properties >>
string path 0.000 27.385 0.000 -0.005 
<< end >>
