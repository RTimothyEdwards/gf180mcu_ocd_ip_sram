magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< psubdiff >>
rect -1382 23 1408 56
rect -1382 -23 -1240 23
rect 1341 -23 1408 23
rect -1382 -56 1408 -23
<< psubdiffcont >>
rect -1240 -23 1341 23
<< metal1 >>
rect -1368 23 1358 41
rect -1368 -23 -1240 23
rect 1341 -23 1358 23
rect -1368 -42 1358 -23
<< end >>
