magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -44 485 44 502
rect -44 -485 -28 485
rect 28 -485 44 485
rect -44 -503 44 -485
<< via2 >>
rect -28 -485 28 485
<< metal3 >>
rect -45 485 45 504
rect -45 -485 -28 485
rect 28 -485 45 485
rect -45 -504 45 -485
<< end >>
