magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< psubdiff >>
rect -55 366 56 400
rect -55 -156 -23 366
rect 23 -156 56 366
rect -55 -190 56 -156
<< psubdiffcont >>
rect -23 -156 23 366
<< metal1 >>
rect -49 366 49 394
rect -49 -156 -23 366
rect 23 -156 49 366
rect -49 -184 49 -156
<< end >>
