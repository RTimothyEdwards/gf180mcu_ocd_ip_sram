magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -1299 104 1299 122
rect -1299 -104 -1283 104
rect 1283 -104 1299 104
rect -1299 -123 1299 -104
<< via2 >>
rect -1283 -104 1283 104
<< metal3 >>
rect -1299 104 1299 123
rect -1299 -104 -1283 104
rect 1283 -104 1299 104
rect -1299 -123 1299 -104
<< end >>
