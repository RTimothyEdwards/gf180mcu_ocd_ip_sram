magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -113 149 113 156
rect -113 -149 -106 149
rect 106 -149 113 149
rect -113 -156 113 -149
<< via2 >>
rect -106 -149 106 149
<< metal3 >>
rect -113 149 113 156
rect -113 -149 -106 149
rect 106 -149 113 149
rect -113 -156 113 -149
<< end >>
