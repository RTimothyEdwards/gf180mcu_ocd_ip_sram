magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal2 >>
rect -107 28 107 46
rect -107 -28 -91 28
rect 91 -28 107 28
rect -107 -46 107 -28
<< via2 >>
rect -91 -28 91 28
<< metal3 >>
rect -108 28 108 46
rect -108 -28 -91 28
rect 91 -28 108 28
rect -108 -46 108 -28
<< end >>
