magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal2 >>
rect -63 28 63 35
rect -63 -28 -56 28
rect 56 -28 63 28
rect -63 -35 63 -28
<< via2 >>
rect -56 -28 56 28
<< metal3 >>
rect -63 28 63 35
rect -63 -28 -56 28
rect 56 -28 63 28
rect -63 -35 63 -28
<< end >>
