magic
tech gf180mcuD
magscale 1 10
timestamp 1764625907
<< metal1 >>
rect 3513 66 3927 122
<< metal3 >>
rect 2538 845 3247 945
rect 2538 635 21443 845
rect 2538 455 3247 635
rect 20927 569 21443 635
rect 2538 -155 3510 335
use M2_M14310591302087_3v1024x8m81  M2_M14310591302087_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2861 0 1 700
box -113 -243 113 243
use M2_M14310591302087_3v1024x8m81  M2_M14310591302087_3v1024x8m81_1
timestamp 1764525316
transform 1 0 3597 0 1 90
box -113 -243 113 243
use M3_M24310591302090_3v1024x8m81  M3_M24310591302090_3v1024x8m81_0
timestamp 1764525316
transform 1 0 3597 0 1 90
box -113 -243 113 243
use M3_M24310591302090_3v1024x8m81  M3_M24310591302090_3v1024x8m81_1
timestamp 1764525316
transform 1 0 2751 0 1 700
box -113 -243 113 243
<< properties >>
string path 25.225 0.500 16.695 0.500 
<< end >>
