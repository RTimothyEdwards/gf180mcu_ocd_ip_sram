magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nwell >>
rect 4608 19539 6692 20186
rect 9694 19994 10581 20197
rect 9694 19940 10808 19994
rect 7130 19545 7550 19596
rect 9695 19550 10808 19940
rect 4608 19504 6273 19539
rect 11564 19517 14760 20166
<< nsubdiff >>
rect 1486 19615 1594 19777
rect 17843 19629 17952 19777
rect 17842 19488 18051 19629
rect 17842 19402 18034 19488
<< polysilicon >>
rect 4589 19864 5251 19920
rect 4589 19788 4661 19864
rect 4485 19760 4661 19788
rect 7730 19780 7969 19788
rect 4485 19732 5251 19760
rect 7730 19732 8050 19780
rect 4592 19704 5251 19732
rect 7879 19724 8050 19732
rect 8358 19724 8451 19780
rect 9564 19745 9637 20043
rect 10754 19780 10826 20082
rect 12782 19864 13445 19920
rect 10713 19724 10826 19780
rect 10908 19725 11108 19780
rect 10908 19724 11028 19725
rect 11423 19724 11928 19781
rect 14707 19780 14779 19921
rect 12782 19704 13445 19760
rect 14707 19724 15356 19780
rect 14707 19704 14779 19724
<< metal1 >>
rect 1486 19675 2811 20070
rect 3026 19850 4435 20121
rect 4537 19770 5359 19854
rect 4537 19727 4618 19770
rect 1404 19615 2811 19675
rect 4368 19643 4618 19727
rect 6521 19727 6602 19943
rect 7969 19828 8339 20107
rect 9471 20013 9828 20107
rect 8404 19829 8919 19877
rect 9456 19829 10160 19877
rect 10687 19809 10961 19855
rect 11028 19805 11398 20107
rect 11659 19968 14659 20052
rect 11659 19839 12581 19968
rect 12788 19727 12849 19896
rect 14628 19789 14828 19836
rect 14926 19815 16342 20107
rect 6521 19643 8339 19727
rect 9499 19670 10170 19716
rect 11028 19643 12849 19727
rect 14746 19696 14828 19789
rect 14746 19650 15411 19696
rect 16625 19688 17952 20070
rect 16625 19615 18034 19688
rect 1404 19358 1506 19615
rect 17932 19401 18034 19615
<< metal2 >>
rect 1464 19403 2947 20147
rect 3885 19403 4442 20094
rect 4515 19403 5416 20094
rect 5730 19403 6346 19732
rect 6713 19403 7130 20094
rect 7193 19403 7658 20094
rect 8075 19403 8292 20094
rect 9795 19655 10181 20094
rect 8428 19365 8847 19508
rect 10518 19403 11120 20107
rect 14078 19403 14919 20094
rect 14994 19403 15565 20107
rect 16484 19403 17973 20147
rect 5992 -14 6083 78
rect 8988 -114 9079 -21
rect 9253 -114 9343 -21
rect 9517 -114 9608 -21
rect 9781 -114 9872 -21
rect 10046 -114 10136 -21
rect 10311 -114 10401 -21
rect 11817 -114 11907 -21
rect 12082 -114 12172 -21
rect 12345 -114 12436 -21
rect 12610 -114 12700 -21
rect 12875 -114 12965 -21
rect 13139 -114 13230 -21
rect 13403 -114 13493 -21
rect 13668 -114 13758 -21
<< metal3 >>
rect 48 19962 139 20055
rect 1443 19928 18161 20069
rect 428 19653 517 19746
rect 1443 19631 3714 19772
rect 5730 19639 9434 19732
rect 48 19362 139 19455
rect 9795 19416 9864 19676
rect 15655 19631 18161 19772
rect 18923 19653 19013 19746
rect 0 19059 89 19152
rect 19348 19059 19438 19152
rect 0 18441 89 18534
rect 19348 18443 19438 18536
rect 0 17847 89 17940
rect 19348 17847 19438 17940
rect 0 17231 89 17324
rect 19348 17231 19438 17324
rect 0 16631 89 16724
rect 19348 16635 19438 16728
rect 0 16015 89 16108
rect 19348 16019 19438 16112
rect 0 15423 89 15516
rect 19348 15423 19438 15516
rect 0 14807 89 14900
rect 19348 14807 19438 14900
rect 0 14211 89 14304
rect 19348 14211 19438 14304
rect 0 13595 89 13688
rect 19348 13595 19438 13688
rect 0 12999 89 13092
rect 19348 12999 19438 13092
rect 0 12383 89 12476
rect 19348 12383 19438 12476
rect 0 11787 89 11880
rect 19348 11787 19438 11880
rect 0 11171 89 11264
rect 19348 11171 19438 11264
rect 0 10575 89 10668
rect 19348 10575 19438 10668
rect 0 9959 89 10052
rect 19348 9959 19438 10052
rect 0 9363 89 9456
rect 19348 9363 19438 9456
rect 0 8747 89 8840
rect 19348 8747 19438 8840
rect 0 8150 89 8243
rect 19348 8151 19438 8244
rect 0 7534 89 7627
rect 19348 7535 19438 7628
rect 0 6939 89 7032
rect 19348 6939 19438 7032
rect 0 6323 89 6416
rect 19348 6323 19438 6416
rect 0 5727 89 5820
rect 19348 5727 19438 5820
rect 0 5111 89 5204
rect 19348 5111 19438 5204
rect 0 4515 89 4608
rect 19348 4515 19438 4608
rect 0 3899 89 3992
rect 19348 3899 19438 3992
rect 0 3301 89 3394
rect 19348 3301 19438 3394
rect 0 2685 89 2778
rect 19348 2685 19438 2778
rect 0 2091 89 2184
rect 19348 2091 19438 2184
rect 0 1475 89 1568
rect 19348 1475 19438 1568
rect 0 880 89 973
rect 19348 881 19438 974
rect 0 263 89 356
rect 19348 265 19438 358
use M1_NACTIVE_02_256x8m81  M1_NACTIVE_02_256x8m81_0
timestamp 1763766357
transform 1 0 9844 0 1 20065
box -54 -56 607 56
use M1_NWELL_01_256x8m81  M1_NWELL_01_256x8m81_0
timestamp 1763766357
transform 1 0 1540 0 1 20014
box -154 -501 1372 159
use M1_NWELL_01_256x8m81  M1_NWELL_01_256x8m81_1
timestamp 1763766357
transform -1 0 17897 0 1 20014
box -154 -501 1372 159
use M1_PACTIVE$10_256x8m81  M1_PACTIVE$10_256x8m81_0
timestamp 1763766357
transform 1 0 8024 0 1 20065
box -54 -56 1271 56
use M1_PACTIVE$10_256x8m81  M1_PACTIVE$10_256x8m81_1
timestamp 1763766357
transform 1 0 3073 0 1 20065
box -54 -56 1271 56
use M1_PACTIVE$10_256x8m81  M1_PACTIVE$10_256x8m81_2
timestamp 1763766357
transform 1 0 15032 0 1 20065
box -54 -56 1271 56
use M1_PACTIVE$11_256x8m81  M1_PACTIVE$11_256x8m81_0
timestamp 1763766357
transform 1 0 11102 0 1 20065
box -54 -56 275 56
use M1_POLY2$$204150828_256x8m81  M1_POLY2$$204150828_256x8m81_0
timestamp 1763766357
transform 1 0 6561 0 1 19812
box -46 -122 46 122
use M1_POLY24310591302019_256x8m81  M1_POLY24310591302019_256x8m81_0
timestamp 1763766357
transform 1 0 8428 0 1 19786
box -36 -80 36 78
use M1_POLY24310591302019_256x8m81  M1_POLY24310591302019_256x8m81_1
timestamp 1763766357
transform 0 -1 9598 1 0 20019
box -36 -80 36 78
use M1_POLY24310591302019_256x8m81  M1_POLY24310591302019_256x8m81_2
timestamp 1763766357
transform 1 0 10937 0 1 19814
box -36 -80 36 78
use M1_POLY24310591302019_256x8m81  M1_POLY24310591302019_256x8m81_3
timestamp 1763766357
transform 1 0 12819 0 1 19814
box -36 -80 36 78
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_0
timestamp 1763766357
transform 1 0 10789 0 1 20052
box -36 -36 36 36
use M2_M1$$201262124_256x8m81  M2_M1$$201262124_256x8m81_0
timestamp 1763766357
transform 1 0 9590 0 1 20017
box -119 -46 119 46
use M2_M1$$204138540_256x8m81  M2_M1$$204138540_256x8m81_0
timestamp 1763766357
transform 1 0 7281 0 1 19847
box -45 -46 340 46
use M2_M1$$204138540_256x8m81  M2_M1$$204138540_256x8m81_1
timestamp 1763766357
transform 1 0 9841 0 1 20060
box -45 -46 340 46
use M2_M1$$204139564_256x8m81  M2_M1$$204139564_256x8m81_0
timestamp 1763766357
transform 1 0 8120 0 1 20027
box -45 -198 171 46
use M2_M1$$204140588_256x8m81  M2_M1$$204140588_256x8m81_0
timestamp 1763766357
transform 1 0 8651 0 1 19685
box -45 -46 783 46
use M2_M1$$204141612_256x8m81  M2_M1$$204141612_256x8m81_0
timestamp 1763766357
transform 1 0 10588 0 1 20060
box -45 -46 487 46
use M2_M1$$204141612_256x8m81  M2_M1$$204141612_256x8m81_1
timestamp 1763766357
transform 1 0 14123 0 1 20010
box -45 -46 487 46
use M2_M1$$204141612_256x8m81  M2_M1$$204141612_256x8m81_2
timestamp 1763766357
transform 1 0 14123 0 1 19685
box -45 -46 487 46
use M2_M1$$204220460_256x8m81  M2_M1$$204220460_256x8m81_0
timestamp 1763766357
transform 1 0 3079 0 1 19687
box -45 -46 635 46
use M2_M1$$204220460_256x8m81  M2_M1$$204220460_256x8m81_1
timestamp 1763766357
transform 1 0 4754 0 1 19975
box -45 -46 635 46
use M2_M1$$204220460_256x8m81  M2_M1$$204220460_256x8m81_2
timestamp 1763766357
transform 1 0 4754 0 1 19650
box -45 -46 635 46
use M2_M1$$204220460_256x8m81  M2_M1$$204220460_256x8m81_3
timestamp 1763766357
transform 1 0 15701 0 1 19685
box -45 -46 635 46
use M2_M1$$204221484_256x8m81  M2_M1$$204221484_256x8m81_0
timestamp 1763766357
transform 1 0 1509 0 1 20024
box -45 -351 1225 46
use M2_M1$$204221484_256x8m81  M2_M1$$204221484_256x8m81_1
timestamp 1763766357
transform -1 0 17928 0 1 20024
box -45 -351 1225 46
use M2_M1$$204222508_256x8m81  M2_M1$$204222508_256x8m81_0
timestamp 1763766357
transform 1 0 3947 0 1 20024
box -45 -198 487 46
use M2_M1$$204222508_256x8m81  M2_M1$$204222508_256x8m81_1
timestamp 1763766357
transform 1 0 15040 0 1 20024
box -45 -198 487 46
use M3_M2$$204142636_256x8m81  M3_M2$$204142636_256x8m81_0
timestamp 1763766357
transform 1 0 3947 0 1 20024
box -44 -46 487 46
use M3_M2$$204142636_256x8m81  M3_M2$$204142636_256x8m81_1
timestamp 1763766357
transform 1 0 5775 0 1 19685
box -44 -46 487 46
use M3_M2$$204142636_256x8m81  M3_M2$$204142636_256x8m81_2
timestamp 1763766357
transform 1 0 15040 0 1 20024
box -44 -46 487 46
use M3_M2$$204142636_256x8m81  M3_M2$$204142636_256x8m81_3
timestamp 1763766357
transform 1 0 15040 0 1 20024
box -44 -46 487 46
use M3_M2$$204143660_256x8m81  M3_M2$$204143660_256x8m81_0
timestamp 1763766357
transform 1 0 8120 0 1 20024
box -45 -46 171 46
use M3_M2$$204144684_256x8m81  M3_M2$$204144684_256x8m81_0
timestamp 1763766357
transform 1 0 3079 0 1 19687
box -45 -46 635 46
use M3_M2$$204144684_256x8m81  M3_M2$$204144684_256x8m81_1
timestamp 1763766357
transform 1 0 15701 0 1 19685
box -45 -46 635 46
use M3_M2$$204145708_256x8m81  M3_M2$$204145708_256x8m81_0
timestamp 1763766357
transform 1 0 8651 0 1 19685
box -45 -46 783 46
use M3_M2$$204146732_256x8m81  M3_M2$$204146732_256x8m81_0
timestamp 1763766357
transform 1 0 9841 0 1 19681
box -45 -46 340 46
use M3_M2$$204147756_256x8m81  M3_M2$$204147756_256x8m81_0
timestamp 1763766357
transform 1 0 8637 0 1 19394
box -193 -46 193 46
use nmos_1p2_01_R270_256x8m81  nmos_1p2_01_R270_256x8m81_0
timestamp 1763766357
transform 0 -1 9522 -1 0 19787
box -102 -44 130 659
use nmos_1p2_02_R90_256x8m81  nmos_1p2_02_R90_256x8m81_0
timestamp 1763766357
transform 0 -1 4442 1 0 19746
box -102 -44 130 987
use nmos_5p04310591302099_256x8m81  nmos_5p04310591302099_256x8m81_0
timestamp 1763766357
transform 0 -1 16342 1 0 19724
box -88 -44 144 987
use nmos_5p043105913020111_256x8m81  nmos_5p043105913020111_256x8m81_0
timestamp 1763766357
transform 0 -1 8339 1 0 19724
box -88 -44 144 291
use nmos_5p043105913020111_256x8m81  nmos_5p043105913020111_256x8m81_1
timestamp 1763766357
transform 0 -1 11398 1 0 19724
box -88 -44 144 291
use pmos_1p2_01_R90_256x8m81  pmos_1p2_01_R90_256x8m81_0
timestamp 1763766357
transform 0 -1 7702 1 0 19746
box -188 -86 216 701
use pmos_1p2_02_R90_256x8m81  pmos_1p2_02_R90_256x8m81_0
timestamp 1763766357
transform 0 -1 6471 1 0 19746
box -216 -86 348 1264
use pmos_1p2_02_R90_256x8m81  pmos_1p2_02_R90_256x8m81_1
timestamp 1763766357
transform 0 -1 14665 1 0 19746
box -216 -86 348 1264
use pmos_5p043105913020101_256x8m81  pmos_5p043105913020101_256x8m81_0
timestamp 1763766357
transform 0 -1 12581 1 0 19724
box -174 -86 230 701
use pmos_5p043105913020101_256x8m81  pmos_5p043105913020101_256x8m81_1
timestamp 1763766357
transform 0 -1 10712 1 0 19724
box -174 -86 230 701
use pmoscap_L1_W2_R270_256x8m81  pmoscap_L1_W2_R270_256x8m81_0
timestamp 1763766357
transform 0 -1 1542 -1 0 20054
box -78 -189 771 1517
use pmoscap_L1_W2_R270_256x8m81  pmoscap_L1_W2_R270_256x8m81_1
timestamp 1763766357
transform 0 1 17896 -1 0 20054
box -78 -189 771 1517
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_0
timestamp 1763766357
transform 0 1 17896 -1 0 10822
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_1
timestamp 1763766357
transform 0 1 17896 -1 0 9610
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_2
timestamp 1763766357
transform 0 1 17896 -1 0 8398
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_3
timestamp 1763766357
transform 0 1 17896 -1 0 7186
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_4
timestamp 1763766357
transform 0 1 17896 -1 0 5974
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_5
timestamp 1763766357
transform 0 1 17896 -1 0 4762
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_6
timestamp 1763766357
transform 0 1 17896 -1 0 3550
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_7
timestamp 1763766357
transform 0 1 17896 -1 0 2338
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_8
timestamp 1763766357
transform 0 1 17896 -1 0 1126
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_9
timestamp 1763766357
transform 0 1 17896 -1 0 19306
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_10
timestamp 1763766357
transform 0 1 17896 -1 0 18094
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_11
timestamp 1763766357
transform 0 1 17896 -1 0 16882
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_12
timestamp 1763766357
transform 0 1 17896 -1 0 15670
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_13
timestamp 1763766357
transform 0 1 17896 -1 0 14458
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_14
timestamp 1763766357
transform 0 1 17896 -1 0 13246
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_15
timestamp 1763766357
transform 0 1 17896 -1 0 12034
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_16
timestamp 1763766357
transform 0 -1 1542 -1 0 10822
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_17
timestamp 1763766357
transform 0 -1 1542 -1 0 9610
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_18
timestamp 1763766357
transform 0 -1 1542 -1 0 8398
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_19
timestamp 1763766357
transform 0 -1 1542 -1 0 7186
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_20
timestamp 1763766357
transform 0 -1 1542 -1 0 5974
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_21
timestamp 1763766357
transform 0 -1 1542 -1 0 4762
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_22
timestamp 1763766357
transform 0 -1 1542 -1 0 3550
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_23
timestamp 1763766357
transform 0 -1 1542 -1 0 2338
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_24
timestamp 1763766357
transform 0 -1 1542 -1 0 1126
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_25
timestamp 1763766357
transform 0 -1 1542 -1 0 19306
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_26
timestamp 1763766357
transform 0 -1 1542 -1 0 18094
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_27
timestamp 1763766357
transform 0 -1 1542 -1 0 16882
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_28
timestamp 1763766357
transform 0 -1 1542 -1 0 15670
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_29
timestamp 1763766357
transform 0 -1 1542 -1 0 14458
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_30
timestamp 1763766357
transform 0 -1 1542 -1 0 13246
box -226 -219 1235 3808
use pmoscap_R270_256x8m81  pmoscap_R270_256x8m81_31
timestamp 1763766357
transform 0 -1 1542 -1 0 12034
box -226 -219 1235 3808
use xdec32_256x8m81  xdec32_256x8m81_0
timestamp 1763766357
transform 1 0 1208 0 1 0
box 230 -159 16952 19575
<< labels >>
rlabel metal2 s 10355 -67 10355 -67 4 xb[0]
port 133 nsew
rlabel metal2 s 10091 -67 10091 -67 4 xb[1]
port 134 nsew
rlabel metal2 s 9827 -67 9827 -67 4 xb[2]
port 135 nsew
rlabel metal2 s 9562 -67 9562 -67 4 xb[3]
port 136 nsew
rlabel metal2 s 11862 -67 11862 -67 4 xa[7]
port 137 nsew
rlabel metal2 s 12126 -67 12126 -67 4 xa[6]
port 138 nsew
rlabel metal2 s 12391 -67 12391 -67 4 xa[5]
port 139 nsew
rlabel metal2 s 12656 -67 12656 -67 4 xa[4]
port 140 nsew
rlabel metal2 s 13713 -67 13713 -67 4 xa[0]
port 141 nsew
rlabel metal2 s 6038 31 6038 31 4 men
port 142 nsew
rlabel metal2 s 12919 -67 12919 -67 4 xa[3]
port 143 nsew
rlabel metal2 s 13184 -67 13184 -67 4 xa[2]
port 144 nsew
rlabel metal2 s 13449 -67 13449 -67 4 xa[1]
port 145 nsew
rlabel metal2 s 9298 -67 9298 -67 4 xc[0]
port 146 nsew
rlabel metal2 s 9034 -67 9034 -67 4 xc[1]
port 147 nsew
rlabel metal3 s 44 927 44 927 4 LWL[1]
port 91 nsew
rlabel metal3 s 44 310 44 310 4 LWL[0]
port 92 nsew
rlabel metal3 s 44 1522 44 1522 4 LWL[2]
port 90 nsew
rlabel metal3 s 44 2138 44 2138 4 LWL[3]
port 89 nsew
rlabel metal3 s 44 2732 44 2732 4 LWL[4]
port 88 nsew
rlabel metal3 s 44 3348 44 3348 4 LWL[5]
port 87 nsew
rlabel metal3 s 44 3946 44 3946 4 LWL[6]
port 95 nsew
rlabel metal3 s 44 4562 44 4562 4 LWL[7]
port 97 nsew
rlabel metal3 s 44 5158 44 5158 4 LWL[8]
port 93 nsew
rlabel metal3 s 44 5774 44 5774 4 LWL[9]
port 94 nsew
rlabel metal3 s 44 6370 44 6370 4 LWL[10]
port 78 nsew
rlabel metal3 s 44 6986 44 6986 4 LWL[11]
port 79 nsew
rlabel metal3 s 44 7581 44 7581 4 LWL[12]
port 80 nsew
rlabel metal3 s 44 8197 44 8197 4 LWL[13]
port 81 nsew
rlabel metal3 s 44 8794 44 8794 4 LWL[14]
port 82 nsew
rlabel metal3 s 44 9410 44 9410 4 LWL[15]
port 83 nsew
rlabel metal3 s 44 10006 44 10006 4 LWL[16]
port 84 nsew
rlabel metal3 s 44 10622 44 10622 4 LWL[17]
port 85 nsew
rlabel metal3 s 44 11218 44 11218 4 LWL[18]
port 86 nsew
rlabel metal3 s 44 11834 44 11834 4 LWL[19]
port 68 nsew
rlabel metal3 s 44 13046 44 13046 4 LWL[21]
port 70 nsew
rlabel metal3 s 44 12430 44 12430 4 LWL[20]
port 69 nsew
rlabel metal3 s 44 13642 44 13642 4 LWL[22]
port 71 nsew
rlabel metal3 s 44 14258 44 14258 4 LWL[23]
port 72 nsew
rlabel metal3 s 44 14854 44 14854 4 LWL[24]
port 73 nsew
rlabel metal3 s 44 15470 44 15470 4 LWL[25]
port 74 nsew
rlabel metal3 s 44 16062 44 16062 4 LWL[26]
port 75 nsew
rlabel metal3 s 44 16678 44 16678 4 LWL[27]
port 76 nsew
rlabel metal3 s 44 18488 44 18488 4 LWL[30]
port 99 nsew
rlabel metal3 s 44 17894 44 17894 4 LWL[29]
port 98 nsew
rlabel metal3 s 44 17278 44 17278 4 LWL[28]
port 77 nsew
rlabel metal3 s 44 19106 44 19106 4 LWL[31]
port 67 nsew
rlabel metal3 s 19393 928 19393 928 4 RWL[1]
port 116 nsew
rlabel metal3 s 19393 312 19393 312 4 RWL[0]
port 115 nsew
rlabel metal3 s 19393 1522 19393 1522 4 RWL[2]
port 114 nsew
rlabel metal3 s 19393 2138 19393 2138 4 RWL[3]
port 117 nsew
rlabel metal3 s 19393 2732 19393 2732 4 RWL[4]
port 113 nsew
rlabel metal3 s 19393 3348 19393 3348 4 RWL[5]
port 118 nsew
rlabel metal3 s 19393 3946 19393 3946 4 RWL[6]
port 112 nsew
rlabel metal3 s 19393 4562 19393 4562 4 RWL[7]
port 119 nsew
rlabel metal3 s 19393 5158 19393 5158 4 RWL[8]
port 120 nsew
rlabel metal3 s 19393 5774 19393 5774 4 RWL[9]
port 121 nsew
rlabel metal3 s 19393 6370 19393 6370 4 RWL[10]
port 122 nsew
rlabel metal3 s 19393 6986 19393 6986 4 RWL[11]
port 123 nsew
rlabel metal3 s 19393 7582 19393 7582 4 RWL[12]
port 124 nsew
rlabel metal3 s 19393 8198 19393 8198 4 RWL[13]
port 125 nsew
rlabel metal3 s 19393 8794 19393 8794 4 RWL[14]
port 126 nsew
rlabel metal3 s 19393 9410 19393 9410 4 RWL[15]
port 127 nsew
rlabel metal3 s 19393 10006 19393 10006 4 RWL[16]
port 128 nsew
rlabel metal3 s 19393 10622 19393 10622 4 RWL[17]
port 129 nsew
rlabel metal3 s 19393 11218 19393 11218 4 RWL[18]
port 130 nsew
rlabel metal3 s 19393 11834 19393 11834 4 RWL[19]
port 131 nsew
rlabel metal3 s 19393 13046 19393 13046 4 RWL[21]
port 111 nsew
rlabel metal3 s 19393 12430 19393 12430 4 RWL[20]
port 132 nsew
rlabel metal3 s 19393 13642 19393 13642 4 RWL[22]
port 110 nsew
rlabel metal3 s 19393 14258 19393 14258 4 RWL[23]
port 109 nsew
rlabel metal3 s 19393 15470 19393 15470 4 RWL[25]
port 107 nsew
rlabel metal3 s 19393 14854 19393 14854 4 RWL[24]
port 108 nsew
rlabel metal3 s 19393 16682 19393 16682 4 RWL[27]
port 105 nsew
rlabel metal3 s 19393 16066 19393 16066 4 RWL[26]
port 106 nsew
rlabel metal3 s 19393 17894 19393 17894 4 RWL[29]
port 103 nsew
rlabel metal3 s 19393 17278 19393 17278 4 RWL[28]
port 104 nsew
rlabel metal3 s 19393 19106 19393 19106 4 RWL[31]
port 101 nsew
rlabel metal3 s 19393 18490 19393 18490 4 RWL[30]
port 102 nsew
rlabel metal3 s 93 20009 93 20009 4 vss
port 64 nsew
rlabel metal3 s 18968 19700 18968 19700 4 DRWL
port 1 nsew
rlabel metal3 s 472 19700 472 19700 4 DLWL
port 66 nsew
rlabel metal3 s 93 19409 93 19409 4 vdd
port 65 nsew
<< end >>
