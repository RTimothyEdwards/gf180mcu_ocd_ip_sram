magic
tech gf180mcuD
magscale 1 10
timestamp 1765833452
<< metal3 >>
rect -1397 19938 -26 19939
rect 124 19938 16315 19939
rect -1397 19687 16315 19938
rect -26 19686 124 19687
rect -1397 19440 -26 19441
rect 124 19440 16315 19441
rect -1397 19189 16315 19440
rect -26 19188 124 19189
rect -1397 18726 -26 18727
rect 124 18726 16315 18727
rect -1397 18475 16315 18726
rect -26 18474 124 18475
rect -1397 18228 -26 18229
rect 124 18228 16315 18229
rect -1397 17977 16315 18228
rect -26 17976 124 17977
rect -1397 17514 -26 17515
rect 124 17514 16315 17515
rect -1397 17263 16315 17514
rect -26 17262 124 17263
rect -1397 17016 -26 17017
rect 124 17016 16315 17017
rect -1397 16765 16315 17016
rect -26 16764 124 16765
rect -1397 16302 -26 16303
rect 124 16302 16315 16303
rect -1397 16051 16315 16302
rect -26 16050 124 16051
rect -1397 15804 -26 15805
rect 124 15804 16315 15805
rect -1397 15553 16315 15804
rect -26 15552 124 15553
rect -1397 15090 -26 15091
rect 124 15090 16315 15091
rect -1397 14839 16315 15090
rect -26 14838 124 14839
rect -1397 14592 -26 14593
rect 124 14592 16315 14593
rect -1397 14341 16315 14592
rect -26 14340 124 14341
rect -1397 13878 -26 13879
rect 124 13878 16315 13879
rect -1397 13627 16315 13878
rect -26 13626 124 13627
rect -1397 13380 -26 13381
rect 124 13380 16315 13381
rect -1397 13129 16315 13380
rect -26 13128 124 13129
rect -1397 12666 -26 12667
rect 124 12666 16315 12667
rect -1397 12415 16315 12666
rect -26 12414 124 12415
rect -1397 12168 -26 12169
rect 124 12168 16315 12169
rect -1397 11917 16315 12168
rect -26 11916 124 11917
rect -1397 11454 -26 11455
rect 124 11454 16315 11455
rect -1397 11203 16315 11454
rect -26 11202 124 11203
rect -1397 10956 -26 10957
rect 124 10956 16315 10957
rect -1397 10705 16315 10956
rect -26 10704 124 10705
rect -1397 10242 -26 10243
rect 124 10242 16315 10243
rect -1397 9991 16315 10242
rect -26 9990 124 9991
rect -1397 9744 -26 9745
rect 124 9744 16315 9745
rect -1397 9493 16315 9744
rect -26 9492 124 9493
rect -1397 9030 -26 9031
rect 124 9030 16315 9031
rect -1397 8779 16315 9030
rect -26 8778 124 8779
rect -1397 8532 -26 8533
rect 124 8532 16315 8533
rect -1397 8281 16315 8532
rect -26 8280 124 8281
rect -1397 7818 -26 7819
rect 124 7818 16315 7819
rect -1397 7567 16315 7818
rect -26 7566 124 7567
rect -1397 7320 -26 7321
rect 124 7320 16315 7321
rect -1397 7069 16315 7320
rect -26 7068 124 7069
rect -1397 6606 -26 6607
rect 124 6606 16315 6607
rect -1397 6355 16315 6606
rect -26 6354 124 6355
rect -1397 6108 -26 6109
rect 124 6108 16315 6109
rect -1397 5857 16315 6108
rect -26 5856 124 5857
rect -1397 5394 -26 5395
rect 124 5394 16315 5395
rect -1397 5143 16315 5394
rect -26 5142 124 5143
rect -1397 4896 -26 4897
rect 124 4896 16315 4897
rect -1397 4645 16315 4896
rect -26 4644 124 4645
rect -1397 4182 -26 4183
rect 124 4182 16315 4183
rect -1397 3931 16315 4182
rect -26 3930 124 3931
rect -1397 3684 -26 3685
rect 124 3684 16315 3685
rect -1397 3433 16315 3684
rect -26 3432 124 3433
rect -1397 2970 -26 2971
rect 124 2970 16315 2971
rect -1397 2719 16315 2970
rect -26 2718 124 2719
rect -1397 2472 -26 2473
rect 124 2472 16315 2473
rect -1397 2221 16315 2472
rect -26 2220 124 2221
rect -1397 1758 -26 1759
rect 124 1758 16315 1759
rect -1397 1507 16315 1758
rect -26 1506 124 1507
rect -1397 1260 -26 1261
rect 124 1260 16315 1261
rect -1397 1009 16315 1260
rect -26 1008 124 1009
rect -1397 247 16315 499
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_0
timestamp 1765833452
transform -1 0 13007 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_1
timestamp 1765833452
transform -1 0 13007 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_2
timestamp 1765833452
transform -1 0 13007 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_3
timestamp 1765833452
transform -1 0 12571 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_4
timestamp 1765833452
transform -1 0 12571 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_5
timestamp 1765833452
transform -1 0 12571 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_6
timestamp 1765833452
transform -1 0 13007 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_7
timestamp 1765833452
transform -1 0 12571 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_8
timestamp 1765833452
transform -1 0 15623 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_9
timestamp 1765833452
transform -1 0 12571 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_10
timestamp 1765833452
transform -1 0 15623 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_11
timestamp 1765833452
transform -1 0 15623 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_12
timestamp 1765833452
transform -1 0 15623 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_13
timestamp 1765833452
transform -1 0 15623 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_14
timestamp 1765833452
transform -1 0 15623 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_15
timestamp 1765833452
transform -1 0 15623 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_16
timestamp 1765833452
transform -1 0 13443 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_17
timestamp 1765833452
transform -1 0 13879 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_18
timestamp 1765833452
transform -1 0 13879 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_19
timestamp 1765833452
transform -1 0 13879 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_20
timestamp 1765833452
transform -1 0 13879 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_21
timestamp 1765833452
transform -1 0 13879 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_22
timestamp 1765833452
transform -1 0 13879 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_23
timestamp 1765833452
transform -1 0 13879 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_24
timestamp 1765833452
transform -1 0 13443 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_25
timestamp 1765833452
transform -1 0 13007 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_26
timestamp 1765833452
transform -1 0 13443 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_27
timestamp 1765833452
transform -1 0 13007 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_28
timestamp 1765833452
transform -1 0 13443 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_29
timestamp 1765833452
transform -1 0 13443 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_30
timestamp 1765833452
transform -1 0 12571 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_31
timestamp 1765833452
transform -1 0 12571 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_32
timestamp 1765833452
transform -1 0 13443 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_33
timestamp 1765833452
transform -1 0 13443 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_34
timestamp 1765833452
transform -1 0 14751 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_35
timestamp 1765833452
transform -1 0 14751 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_36
timestamp 1765833452
transform -1 0 14315 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_37
timestamp 1765833452
transform -1 0 14315 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_38
timestamp 1765833452
transform -1 0 14315 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_39
timestamp 1765833452
transform -1 0 14315 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_40
timestamp 1765833452
transform -1 0 15187 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_41
timestamp 1765833452
transform -1 0 15187 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_42
timestamp 1765833452
transform -1 0 15187 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_43
timestamp 1765833452
transform -1 0 15187 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_44
timestamp 1765833452
transform -1 0 15187 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_45
timestamp 1765833452
transform -1 0 15187 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_46
timestamp 1765833452
transform -1 0 15187 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_47
timestamp 1765833452
transform -1 0 14315 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_48
timestamp 1765833452
transform -1 0 14315 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_49
timestamp 1765833452
transform -1 0 14315 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_50
timestamp 1765833452
transform -1 0 13007 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_51
timestamp 1765833452
transform -1 0 14751 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_52
timestamp 1765833452
transform -1 0 14751 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_53
timestamp 1765833452
transform -1 0 14751 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_54
timestamp 1765833452
transform -1 0 14751 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_55
timestamp 1765833452
transform -1 0 14751 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_56
timestamp 1765833452
transform 1 0 8063 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_57
timestamp 1765833452
transform 1 0 8063 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_58
timestamp 1765833452
transform 1 0 8063 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_59
timestamp 1765833452
transform 1 0 8063 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_60
timestamp 1765833452
transform 1 0 8063 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_61
timestamp 1765833452
transform 1 0 8063 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_62
timestamp 1765833452
transform 1 0 8063 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_63
timestamp 1765833452
transform 1 0 8499 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_64
timestamp 1765833452
transform 1 0 8499 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_65
timestamp 1765833452
transform 1 0 8499 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_66
timestamp 1765833452
transform 1 0 10679 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_67
timestamp 1765833452
transform 1 0 10243 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_68
timestamp 1765833452
transform 1 0 10679 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_69
timestamp 1765833452
transform 1 0 10679 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_70
timestamp 1765833452
transform 1 0 10679 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_71
timestamp 1765833452
transform 1 0 10679 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_72
timestamp 1765833452
transform 1 0 8935 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_73
timestamp 1765833452
transform 1 0 8935 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_74
timestamp 1765833452
transform 1 0 8935 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_75
timestamp 1765833452
transform 1 0 8935 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_76
timestamp 1765833452
transform 1 0 10243 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_77
timestamp 1765833452
transform 1 0 10243 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_78
timestamp 1765833452
transform 1 0 10243 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_79
timestamp 1765833452
transform 1 0 10243 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_80
timestamp 1765833452
transform 1 0 10243 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_81
timestamp 1765833452
transform 1 0 10243 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_82
timestamp 1765833452
transform 1 0 8935 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_83
timestamp 1765833452
transform 1 0 10679 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_84
timestamp 1765833452
transform 1 0 9807 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_85
timestamp 1765833452
transform 1 0 9807 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_86
timestamp 1765833452
transform 1 0 9807 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_87
timestamp 1765833452
transform 1 0 9807 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_88
timestamp 1765833452
transform 1 0 9807 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_89
timestamp 1765833452
transform 1 0 10679 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_90
timestamp 1765833452
transform 1 0 11115 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_91
timestamp 1765833452
transform 1 0 11115 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_92
timestamp 1765833452
transform 1 0 11115 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_93
timestamp 1765833452
transform 1 0 11115 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_94
timestamp 1765833452
transform 1 0 11115 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_95
timestamp 1765833452
transform 1 0 11115 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_96
timestamp 1765833452
transform 1 0 11115 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_97
timestamp 1765833452
transform 1 0 9807 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_98
timestamp 1765833452
transform 1 0 9807 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_99
timestamp 1765833452
transform 1 0 9371 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_100
timestamp 1765833452
transform 1 0 9371 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_101
timestamp 1765833452
transform 1 0 9371 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_102
timestamp 1765833452
transform 1 0 9371 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_103
timestamp 1765833452
transform 1 0 9371 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_104
timestamp 1765833452
transform 1 0 9371 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_105
timestamp 1765833452
transform 1 0 9371 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_106
timestamp 1765833452
transform 1 0 8499 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_107
timestamp 1765833452
transform 1 0 8499 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_108
timestamp 1765833452
transform 1 0 8499 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_109
timestamp 1765833452
transform 1 0 8499 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_110
timestamp 1765833452
transform 1 0 8935 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_111
timestamp 1765833452
transform 1 0 8935 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_112
timestamp 1765833452
transform 1 0 11115 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_113
timestamp 1765833452
transform 1 0 8063 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_114
timestamp 1765833452
transform 1 0 11115 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_115
timestamp 1765833452
transform 1 0 11115 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_116
timestamp 1765833452
transform 1 0 11115 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_117
timestamp 1765833452
transform 1 0 9371 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_118
timestamp 1765833452
transform 1 0 11115 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_119
timestamp 1765833452
transform 1 0 9371 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_120
timestamp 1765833452
transform 1 0 8063 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_121
timestamp 1765833452
transform 1 0 8063 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_122
timestamp 1765833452
transform 1 0 9371 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_123
timestamp 1765833452
transform 1 0 10679 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_124
timestamp 1765833452
transform 1 0 10679 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_125
timestamp 1765833452
transform 1 0 9371 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_126
timestamp 1765833452
transform 1 0 9371 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_127
timestamp 1765833452
transform 1 0 8499 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_128
timestamp 1765833452
transform 1 0 8499 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_129
timestamp 1765833452
transform 1 0 10679 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_130
timestamp 1765833452
transform 1 0 10679 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_131
timestamp 1765833452
transform 1 0 10679 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_132
timestamp 1765833452
transform 1 0 10679 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_133
timestamp 1765833452
transform 1 0 9371 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_134
timestamp 1765833452
transform 1 0 11115 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_135
timestamp 1765833452
transform 1 0 8499 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_136
timestamp 1765833452
transform 1 0 8935 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_137
timestamp 1765833452
transform 1 0 10243 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_138
timestamp 1765833452
transform 1 0 10243 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_139
timestamp 1765833452
transform 1 0 10243 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_140
timestamp 1765833452
transform 1 0 10243 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_141
timestamp 1765833452
transform 1 0 10243 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_142
timestamp 1765833452
transform 1 0 10243 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_143
timestamp 1765833452
transform 1 0 8063 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_144
timestamp 1765833452
transform 1 0 8063 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_145
timestamp 1765833452
transform 1 0 8935 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_146
timestamp 1765833452
transform 1 0 8935 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_147
timestamp 1765833452
transform 1 0 8935 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_148
timestamp 1765833452
transform 1 0 8935 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_149
timestamp 1765833452
transform 1 0 8935 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_150
timestamp 1765833452
transform 1 0 9807 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_151
timestamp 1765833452
transform 1 0 9807 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_152
timestamp 1765833452
transform 1 0 9807 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_153
timestamp 1765833452
transform 1 0 9807 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_154
timestamp 1765833452
transform 1 0 9807 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_155
timestamp 1765833452
transform 1 0 9807 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_156
timestamp 1765833452
transform 1 0 8499 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_157
timestamp 1765833452
transform 1 0 8499 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_158
timestamp 1765833452
transform 1 0 8499 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_159
timestamp 1765833452
transform 1 0 8063 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_160
timestamp 1765833452
transform -1 0 13007 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_161
timestamp 1765833452
transform -1 0 14751 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_162
timestamp 1765833452
transform -1 0 13007 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_163
timestamp 1765833452
transform -1 0 13007 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_164
timestamp 1765833452
transform -1 0 13007 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_165
timestamp 1765833452
transform -1 0 13007 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_166
timestamp 1765833452
transform -1 0 13007 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_167
timestamp 1765833452
transform -1 0 14751 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_168
timestamp 1765833452
transform -1 0 14315 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_169
timestamp 1765833452
transform -1 0 14315 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_170
timestamp 1765833452
transform -1 0 13443 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_171
timestamp 1765833452
transform -1 0 12571 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_172
timestamp 1765833452
transform -1 0 12571 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_173
timestamp 1765833452
transform -1 0 12571 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_174
timestamp 1765833452
transform -1 0 12571 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_175
timestamp 1765833452
transform -1 0 12571 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_176
timestamp 1765833452
transform -1 0 12571 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_177
timestamp 1765833452
transform -1 0 13443 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_178
timestamp 1765833452
transform -1 0 13443 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_179
timestamp 1765833452
transform -1 0 13443 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_180
timestamp 1765833452
transform -1 0 13443 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_181
timestamp 1765833452
transform -1 0 13443 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_182
timestamp 1765833452
transform -1 0 14315 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_183
timestamp 1765833452
transform -1 0 15623 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_184
timestamp 1765833452
transform -1 0 15623 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_185
timestamp 1765833452
transform -1 0 15623 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_186
timestamp 1765833452
transform -1 0 15623 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_187
timestamp 1765833452
transform -1 0 15623 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_188
timestamp 1765833452
transform -1 0 15623 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_189
timestamp 1765833452
transform -1 0 14315 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_190
timestamp 1765833452
transform -1 0 14315 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_191
timestamp 1765833452
transform -1 0 14315 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_192
timestamp 1765833452
transform -1 0 14751 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_193
timestamp 1765833452
transform -1 0 15187 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_194
timestamp 1765833452
transform -1 0 15187 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_195
timestamp 1765833452
transform -1 0 15187 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_196
timestamp 1765833452
transform -1 0 15187 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_197
timestamp 1765833452
transform -1 0 15187 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_198
timestamp 1765833452
transform -1 0 15187 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_199
timestamp 1765833452
transform -1 0 14751 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_200
timestamp 1765833452
transform -1 0 14751 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_201
timestamp 1765833452
transform -1 0 14751 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_202
timestamp 1765833452
transform -1 0 13879 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_203
timestamp 1765833452
transform -1 0 13879 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_204
timestamp 1765833452
transform -1 0 13879 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_205
timestamp 1765833452
transform -1 0 13879 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_206
timestamp 1765833452
transform -1 0 13879 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_207
timestamp 1765833452
transform -1 0 13879 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_208
timestamp 1765833452
transform -1 0 13007 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_209
timestamp 1765833452
transform -1 0 13007 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_210
timestamp 1765833452
transform -1 0 12571 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_211
timestamp 1765833452
transform -1 0 12571 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_212
timestamp 1765833452
transform 1 0 9807 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_213
timestamp 1765833452
transform 1 0 9807 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_214
timestamp 1765833452
transform 1 0 8063 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_215
timestamp 1765833452
transform 1 0 8063 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_216
timestamp 1765833452
transform -1 0 15623 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_217
timestamp 1765833452
transform -1 0 15623 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_218
timestamp 1765833452
transform 1 0 10243 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_219
timestamp 1765833452
transform 1 0 10243 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_220
timestamp 1765833452
transform -1 0 15187 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_221
timestamp 1765833452
transform -1 0 15187 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_222
timestamp 1765833452
transform -1 0 13879 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_223
timestamp 1765833452
transform -1 0 13879 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_224
timestamp 1765833452
transform 1 0 8935 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_225
timestamp 1765833452
transform 1 0 8935 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_226
timestamp 1765833452
transform -1 0 13443 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_227
timestamp 1765833452
transform -1 0 13443 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_228
timestamp 1765833452
transform 1 0 10679 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_229
timestamp 1765833452
transform 1 0 10679 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_230
timestamp 1765833452
transform -1 0 14751 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_231
timestamp 1765833452
transform -1 0 14751 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_232
timestamp 1765833452
transform 1 0 8499 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_233
timestamp 1765833452
transform 1 0 8499 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_234
timestamp 1765833452
transform -1 0 14315 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_235
timestamp 1765833452
transform -1 0 14315 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_236
timestamp 1765833452
transform 1 0 9371 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_237
timestamp 1765833452
transform 1 0 9371 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_238
timestamp 1765833452
transform 1 0 11115 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_239
timestamp 1765833452
transform 1 0 11115 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_240
timestamp 1765833452
transform -1 0 6935 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_241
timestamp 1765833452
transform -1 0 6935 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_242
timestamp 1765833452
transform -1 0 6935 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_243
timestamp 1765833452
transform -1 0 6935 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_244
timestamp 1765833452
transform -1 0 6935 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_245
timestamp 1765833452
transform -1 0 6935 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_246
timestamp 1765833452
transform -1 0 6935 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_247
timestamp 1765833452
transform -1 0 7807 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_248
timestamp 1765833452
transform -1 0 7807 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_249
timestamp 1765833452
transform -1 0 7807 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_250
timestamp 1765833452
transform -1 0 5627 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_251
timestamp 1765833452
transform -1 0 5627 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_252
timestamp 1765833452
transform -1 0 5627 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_253
timestamp 1765833452
transform -1 0 5627 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_254
timestamp 1765833452
transform -1 0 5627 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_255
timestamp 1765833452
transform -1 0 5627 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_257
timestamp 1765833452
transform -1 0 4755 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_258
timestamp 1765833452
transform -1 0 4755 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_259
timestamp 1765833452
transform -1 0 4755 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_260
timestamp 1765833452
transform -1 0 4755 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_261
timestamp 1765833452
transform -1 0 4755 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_262
timestamp 1765833452
transform -1 0 4755 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_263
timestamp 1765833452
transform -1 0 4755 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_264
timestamp 1765833452
transform -1 0 7807 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_265
timestamp 1765833452
transform -1 0 7807 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_266
timestamp 1765833452
transform -1 0 7807 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_267
timestamp 1765833452
transform -1 0 7807 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_268
timestamp 1765833452
transform -1 0 7371 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_269
timestamp 1765833452
transform -1 0 7371 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_270
timestamp 1765833452
transform -1 0 7371 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_271
timestamp 1765833452
transform -1 0 7371 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_272
timestamp 1765833452
transform -1 0 7371 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_273
timestamp 1765833452
transform -1 0 7371 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_274
timestamp 1765833452
transform -1 0 7371 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_275
timestamp 1765833452
transform -1 0 6063 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_276
timestamp 1765833452
transform -1 0 6063 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_277
timestamp 1765833452
transform -1 0 6063 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_278
timestamp 1765833452
transform -1 0 6499 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_279
timestamp 1765833452
transform -1 0 6499 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_280
timestamp 1765833452
transform -1 0 6499 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_281
timestamp 1765833452
transform -1 0 6499 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_282
timestamp 1765833452
transform -1 0 5191 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_283
timestamp 1765833452
transform -1 0 5191 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_284
timestamp 1765833452
transform -1 0 5191 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_285
timestamp 1765833452
transform -1 0 5191 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_286
timestamp 1765833452
transform -1 0 5191 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_287
timestamp 1765833452
transform -1 0 5191 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_288
timestamp 1765833452
transform -1 0 5191 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_289
timestamp 1765833452
transform -1 0 6499 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_290
timestamp 1765833452
transform -1 0 6499 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_291
timestamp 1765833452
transform -1 0 6499 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_292
timestamp 1765833452
transform -1 0 6063 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_293
timestamp 1765833452
transform -1 0 6063 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_294
timestamp 1765833452
transform -1 0 6063 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_295
timestamp 1765833452
transform -1 0 6063 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_296
timestamp 1765833452
transform 1 0 1119 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_297
timestamp 1765833452
transform 1 0 247 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_298
timestamp 1765833452
transform 1 0 247 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_299
timestamp 1765833452
transform 1 0 247 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_300
timestamp 1765833452
transform 1 0 1555 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_301
timestamp 1765833452
transform 1 0 1555 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_302
timestamp 1765833452
transform 1 0 1555 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_303
timestamp 1765833452
transform 1 0 1555 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_304
timestamp 1765833452
transform 1 0 1555 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_305
timestamp 1765833452
transform 1 0 1555 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_306
timestamp 1765833452
transform 1 0 247 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_307
timestamp 1765833452
transform 1 0 247 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_308
timestamp 1765833452
transform 1 0 247 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_309
timestamp 1765833452
transform 1 0 683 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_310
timestamp 1765833452
transform 1 0 683 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_311
timestamp 1765833452
transform 1 0 683 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_312
timestamp 1765833452
transform 1 0 3299 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_313
timestamp 1765833452
transform 1 0 3299 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_314
timestamp 1765833452
transform 1 0 3299 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_315
timestamp 1765833452
transform 1 0 3299 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_316
timestamp 1765833452
transform 1 0 3299 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_317
timestamp 1765833452
transform 1 0 3299 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_318
timestamp 1765833452
transform 1 0 3299 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_319
timestamp 1765833452
transform 1 0 683 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_320
timestamp 1765833452
transform 1 0 683 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_321
timestamp 1765833452
transform 1 0 2863 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_322
timestamp 1765833452
transform 1 0 2863 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_323
timestamp 1765833452
transform 1 0 2863 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_324
timestamp 1765833452
transform 1 0 2863 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_325
timestamp 1765833452
transform 1 0 2863 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_326
timestamp 1765833452
transform 1 0 683 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_327
timestamp 1765833452
transform 1 0 1991 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_328
timestamp 1765833452
transform 1 0 1991 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_329
timestamp 1765833452
transform 1 0 1991 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_330
timestamp 1765833452
transform 1 0 1991 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_331
timestamp 1765833452
transform 1 0 2863 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_332
timestamp 1765833452
transform 1 0 2863 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_333
timestamp 1765833452
transform 1 0 1991 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_334
timestamp 1765833452
transform 1 0 1991 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_335
timestamp 1765833452
transform 1 0 1991 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_336
timestamp 1765833452
transform 1 0 2427 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_337
timestamp 1765833452
transform 1 0 2427 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_338
timestamp 1765833452
transform 1 0 2427 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_339
timestamp 1765833452
transform 1 0 2427 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_340
timestamp 1765833452
transform 1 0 2427 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_341
timestamp 1765833452
transform 1 0 1555 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_342
timestamp 1765833452
transform 1 0 2427 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_343
timestamp 1765833452
transform 1 0 2427 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_344
timestamp 1765833452
transform 1 0 683 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_345
timestamp 1765833452
transform 1 0 1119 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_346
timestamp 1765833452
transform 1 0 247 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_347
timestamp 1765833452
transform 1 0 1119 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_348
timestamp 1765833452
transform 1 0 1119 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_349
timestamp 1765833452
transform 1 0 1119 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_350
timestamp 1765833452
transform 1 0 1119 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_351
timestamp 1765833452
transform 1 0 1119 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_352
timestamp 1765833452
transform 1 0 683 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_353
timestamp 1765833452
transform 1 0 683 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_354
timestamp 1765833452
transform 1 0 683 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_355
timestamp 1765833452
transform 1 0 3299 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_356
timestamp 1765833452
transform 1 0 3299 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_357
timestamp 1765833452
transform 1 0 3299 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_358
timestamp 1765833452
transform 1 0 3299 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_359
timestamp 1765833452
transform 1 0 3299 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_360
timestamp 1765833452
transform 1 0 1555 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_361
timestamp 1765833452
transform 1 0 1555 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_362
timestamp 1765833452
transform 1 0 1555 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_363
timestamp 1765833452
transform 1 0 1555 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_364
timestamp 1765833452
transform 1 0 1555 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_365
timestamp 1765833452
transform 1 0 1555 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_366
timestamp 1765833452
transform 1 0 2427 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_367
timestamp 1765833452
transform 1 0 2427 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_368
timestamp 1765833452
transform 1 0 2427 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_369
timestamp 1765833452
transform 1 0 2427 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_370
timestamp 1765833452
transform 1 0 2427 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_371
timestamp 1765833452
transform 1 0 683 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_372
timestamp 1765833452
transform 1 0 683 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_373
timestamp 1765833452
transform 1 0 3299 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_374
timestamp 1765833452
transform 1 0 247 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_375
timestamp 1765833452
transform 1 0 247 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_376
timestamp 1765833452
transform 1 0 247 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_377
timestamp 1765833452
transform 1 0 247 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_378
timestamp 1765833452
transform 1 0 2427 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_379
timestamp 1765833452
transform 1 0 1119 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_380
timestamp 1765833452
transform 1 0 2863 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_381
timestamp 1765833452
transform 1 0 2863 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_382
timestamp 1765833452
transform 1 0 2863 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_383
timestamp 1765833452
transform 1 0 2863 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_384
timestamp 1765833452
transform 1 0 2863 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_385
timestamp 1765833452
transform 1 0 2863 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_386
timestamp 1765833452
transform 1 0 1991 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_387
timestamp 1765833452
transform 1 0 1991 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_388
timestamp 1765833452
transform 1 0 1991 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_389
timestamp 1765833452
transform 1 0 1991 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_390
timestamp 1765833452
transform 1 0 1991 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_391
timestamp 1765833452
transform 1 0 1991 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_392
timestamp 1765833452
transform 1 0 247 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_393
timestamp 1765833452
transform 1 0 247 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_394
timestamp 1765833452
transform 1 0 1119 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_395
timestamp 1765833452
transform 1 0 1119 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_396
timestamp 1765833452
transform 1 0 1119 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_397
timestamp 1765833452
transform 1 0 1119 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_398
timestamp 1765833452
transform 1 0 1119 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_399
timestamp 1765833452
transform 1 0 683 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_400
timestamp 1765833452
transform -1 0 7371 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_401
timestamp 1765833452
transform -1 0 7371 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_402
timestamp 1765833452
transform -1 0 7371 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_403
timestamp 1765833452
transform -1 0 7371 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_404
timestamp 1765833452
transform -1 0 7371 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_405
timestamp 1765833452
transform -1 0 7371 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_406
timestamp 1765833452
transform -1 0 7807 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_407
timestamp 1765833452
transform -1 0 7807 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_408
timestamp 1765833452
transform -1 0 7807 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_409
timestamp 1765833452
transform -1 0 6063 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_410
timestamp 1765833452
transform -1 0 6063 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_411
timestamp 1765833452
transform -1 0 5191 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_412
timestamp 1765833452
transform -1 0 5191 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_413
timestamp 1765833452
transform -1 0 5191 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_414
timestamp 1765833452
transform -1 0 5191 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_415
timestamp 1765833452
transform -1 0 5191 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_416
timestamp 1765833452
transform -1 0 5191 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_417
timestamp 1765833452
transform -1 0 6063 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_418
timestamp 1765833452
transform -1 0 6063 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_419
timestamp 1765833452
transform -1 0 6063 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_420
timestamp 1765833452
transform -1 0 6063 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_421
timestamp 1765833452
transform -1 0 4755 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_422
timestamp 1765833452
transform -1 0 4755 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_423
timestamp 1765833452
transform -1 0 4755 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_424
timestamp 1765833452
transform -1 0 4755 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_425
timestamp 1765833452
transform -1 0 4755 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_426
timestamp 1765833452
transform -1 0 4755 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_427
timestamp 1765833452
transform -1 0 7807 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_428
timestamp 1765833452
transform -1 0 7807 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_429
timestamp 1765833452
transform -1 0 7807 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_430
timestamp 1765833452
transform -1 0 5627 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_431
timestamp 1765833452
transform -1 0 6935 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_432
timestamp 1765833452
transform -1 0 6935 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_433
timestamp 1765833452
transform -1 0 6935 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_434
timestamp 1765833452
transform -1 0 6935 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_435
timestamp 1765833452
transform -1 0 6935 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_436
timestamp 1765833452
transform -1 0 6935 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_437
timestamp 1765833452
transform -1 0 5627 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_438
timestamp 1765833452
transform -1 0 5627 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_439
timestamp 1765833452
transform -1 0 5627 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_440
timestamp 1765833452
transform -1 0 5627 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_441
timestamp 1765833452
transform -1 0 6499 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_442
timestamp 1765833452
transform -1 0 6499 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_443
timestamp 1765833452
transform -1 0 6499 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_444
timestamp 1765833452
transform -1 0 6499 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_445
timestamp 1765833452
transform -1 0 6499 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_446
timestamp 1765833452
transform -1 0 6499 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_447
timestamp 1765833452
transform -1 0 5627 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_448
timestamp 1765833452
transform 1 0 1555 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_449
timestamp 1765833452
transform 1 0 1555 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_450
timestamp 1765833452
transform -1 0 5191 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_451
timestamp 1765833452
transform -1 0 5191 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_452
timestamp 1765833452
transform 1 0 2863 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_453
timestamp 1765833452
transform 1 0 2863 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_454
timestamp 1765833452
transform -1 0 4755 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_455
timestamp 1765833452
transform -1 0 4755 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_456
timestamp 1765833452
transform 1 0 247 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_457
timestamp 1765833452
transform 1 0 247 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_458
timestamp 1765833452
transform -1 0 6935 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_459
timestamp 1765833452
transform -1 0 6935 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_460
timestamp 1765833452
transform 1 0 3299 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_461
timestamp 1765833452
transform 1 0 3299 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_462
timestamp 1765833452
transform -1 0 6499 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_463
timestamp 1765833452
transform -1 0 6499 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_464
timestamp 1765833452
transform 1 0 1991 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_465
timestamp 1765833452
transform -1 0 6063 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_466
timestamp 1765833452
transform -1 0 6063 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_467
timestamp 1765833452
transform 1 0 1991 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_468
timestamp 1765833452
transform -1 0 5627 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_469
timestamp 1765833452
transform -1 0 5627 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_470
timestamp 1765833452
transform 1 0 1119 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_471
timestamp 1765833452
transform 1 0 1119 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_472
timestamp 1765833452
transform 1 0 683 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_473
timestamp 1765833452
transform -1 0 7807 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_474
timestamp 1765833452
transform -1 0 7807 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_475
timestamp 1765833452
transform 1 0 683 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_476
timestamp 1765833452
transform 1 0 2427 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_477
timestamp 1765833452
transform 1 0 2427 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_478
timestamp 1765833452
transform -1 0 7371 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_479
timestamp 1765833452
transform -1 0 7371 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_512
timestamp 1765833452
transform -1 0 5627 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_960
timestamp 1765833452
transform -1 0 13007 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_962
timestamp 1765833452
transform -1 0 12571 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_964
timestamp 1765833452
transform -1 0 5191 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_966
timestamp 1765833452
transform -1 0 4755 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_968
timestamp 1765833452
transform -1 0 6935 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_970
timestamp 1765833452
transform -1 0 6499 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_972
timestamp 1765833452
transform -1 0 6063 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_974
timestamp 1765833452
transform -1 0 5627 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_976
timestamp 1765833452
transform -1 0 7807 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_978
timestamp 1765833452
transform -1 0 7371 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_980
timestamp 1765833452
transform -1 0 15623 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_982
timestamp 1765833452
transform -1 0 15187 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_984
timestamp 1765833452
transform -1 0 13879 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_986
timestamp 1765833452
transform -1 0 13443 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_988
timestamp 1765833452
transform -1 0 14751 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_990
timestamp 1765833452
transform -1 0 14315 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_992
timestamp 1765833452
transform 1 0 1119 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_994
timestamp 1765833452
transform 1 0 1555 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_996
timestamp 1765833452
transform 1 0 2863 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_998
timestamp 1765833452
transform 1 0 3299 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_1000
timestamp 1765833452
transform 1 0 1991 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_1002
timestamp 1765833452
transform 1 0 2427 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_1004
timestamp 1765833452
transform 1 0 247 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_1006
timestamp 1765833452
transform 1 0 683 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_1008
timestamp 1765833452
transform 1 0 10679 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_1010
timestamp 1765833452
transform 1 0 11115 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_1012
timestamp 1765833452
transform 1 0 9807 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_1014
timestamp 1765833452
transform 1 0 10243 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_1016
timestamp 1765833452
transform 1 0 8935 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_1018
timestamp 1765833452
transform 1 0 9371 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_1020
timestamp 1765833452
transform 1 0 8063 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v256x8m81  018SRAM_cell1_2x_3v256x8m81_1022
timestamp 1765833452
transform 1 0 8499 0 1 18180
box 30 103 570 1445
use 018SRAM_strap1_2x_3v256x8m81  018SRAM_strap1_2x_3v256x8m81_0
array 0 0 -420 0 15 1212
timestamp 1765833452
transform -1 0 8236 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_2x_3v256x8m81  018SRAM_strap1_2x_3v256x8m81_1
array 0 0 -420 0 15 1212
timestamp 1765833452
transform -1 0 12144 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_2x_3v256x8m81  018SRAM_strap1_2x_3v256x8m81_3
array 0 0 -420 0 15 1212
timestamp 1765833452
transform -1 0 4328 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_0
timestamp 1765833244
transform 1 0 15450 0 1 6708
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_1
timestamp 1765833244
transform 1 0 15450 0 -1 9384
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_2
timestamp 1765833244
transform 1 0 15450 0 -1 8172
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_3
timestamp 1765833244
transform 1 0 15450 0 -1 6960
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_4
timestamp 1765833244
transform 1 0 15450 0 -1 5748
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_5
timestamp 1765833244
transform 1 0 15450 0 -1 4536
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_6
timestamp 1765833244
transform 1 0 15450 0 -1 3324
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_7
timestamp 1765833244
transform 1 0 15450 0 -1 2112
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_8
timestamp 1765833244
transform 1 0 15450 0 -1 900
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_9
timestamp 1765833244
transform 1 0 15450 0 1 648
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_10
timestamp 1765833244
transform 1 0 15450 0 1 1860
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_11
timestamp 1765833244
transform 1 0 15450 0 1 3072
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_12
timestamp 1765833244
transform 1 0 15450 0 1 4284
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_13
timestamp 1765833244
transform 1 0 15450 0 1 7920
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_14
timestamp 1765833244
transform 1 0 15450 0 1 5496
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_15
timestamp 1765833244
transform 1 0 15450 0 1 10344
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_16
timestamp 1765833244
transform 1 0 15450 0 1 11556
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_17
timestamp 1765833244
transform 1 0 15450 0 1 12768
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_18
timestamp 1765833244
transform 1 0 15450 0 1 13980
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_19
timestamp 1765833244
transform 1 0 15450 0 1 15192
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_20
timestamp 1765833244
transform 1 0 15450 0 1 16404
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_21
timestamp 1765833244
transform 1 0 15450 0 1 17616
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_22
timestamp 1765833244
transform 1 0 15450 0 -1 19080
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_23
timestamp 1765833244
transform 1 0 15450 0 -1 17868
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_24
timestamp 1765833244
transform 1 0 15450 0 -1 16656
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_25
timestamp 1765833244
transform 1 0 15450 0 -1 15444
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_26
timestamp 1765833244
transform 1 0 15450 0 -1 14232
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_27
timestamp 1765833244
transform 1 0 15450 0 -1 13020
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_28
timestamp 1765833244
transform 1 0 15450 0 -1 11808
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_29
timestamp 1765833244
transform 1 0 15450 0 1 9132
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_30
timestamp 1765833244
transform 1 0 15450 0 -1 10596
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_31
timestamp 1765833244
transform -1 0 420 0 -1 5748
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_32
timestamp 1765833244
transform -1 0 420 0 -1 4536
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_33
timestamp 1765833244
transform -1 0 420 0 -1 3324
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_34
timestamp 1765833244
transform -1 0 420 0 -1 2112
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_35
timestamp 1765833244
transform -1 0 420 0 -1 900
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_36
timestamp 1765833244
transform -1 0 420 0 1 648
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_37
timestamp 1765833244
transform -1 0 420 0 1 1860
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_38
timestamp 1765833244
transform -1 0 420 0 1 3072
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_39
timestamp 1765833244
transform -1 0 420 0 1 4284
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_40
timestamp 1765833244
transform -1 0 420 0 1 5496
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_41
timestamp 1765833244
transform -1 0 420 0 1 6708
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_42
timestamp 1765833244
transform -1 0 420 0 1 7920
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_43
timestamp 1765833244
transform -1 0 420 0 -1 9384
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_44
timestamp 1765833244
transform -1 0 420 0 -1 8172
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_45
timestamp 1765833244
transform -1 0 420 0 -1 6960
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_46
timestamp 1765833244
transform -1 0 420 0 1 16404
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_47
timestamp 1765833244
transform -1 0 420 0 1 17616
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_48
timestamp 1765833244
transform -1 0 420 0 -1 19080
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_49
timestamp 1765833244
transform -1 0 420 0 -1 17868
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_50
timestamp 1765833244
transform -1 0 420 0 1 10344
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_51
timestamp 1765833244
transform -1 0 420 0 1 11556
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_52
timestamp 1765833244
transform -1 0 420 0 1 12768
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_53
timestamp 1765833244
transform -1 0 420 0 1 13980
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_54
timestamp 1765833244
transform -1 0 420 0 1 15192
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_55
timestamp 1765833244
transform -1 0 420 0 -1 16656
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_56
timestamp 1765833244
transform -1 0 420 0 -1 15444
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_57
timestamp 1765833244
transform -1 0 420 0 -1 14232
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_58
timestamp 1765833244
transform -1 0 420 0 -1 13020
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_59
timestamp 1765833244
transform -1 0 420 0 -1 11808
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_60
timestamp 1765833244
transform -1 0 420 0 1 9132
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_61
timestamp 1765833244
transform -1 0 420 0 -1 10596
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_124
timestamp 1765833244
transform -1 0 420 0 1 18828
box 91 55 511 797
use 018SRAM_strap1_bndry_3v256x8m81  018SRAM_strap1_bndry_3v256x8m81_127
timestamp 1765833244
transform 1 0 15450 0 1 18828
box 91 55 511 797
<< end >>
