magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< nwell >>
rect -133 -66 160 1335
<< polysilicon >>
rect -14 1269 41 1303
rect -14 -34 41 0
use pmos_5p0431059130204_3v512x8m81  pmos_5p0431059130204_3v512x8m81_0
timestamp 1764525316
transform 1 0 -14 0 1 0
box -174 -86 230 1356
<< end >>
