magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -44 104 44 122
rect -44 -104 -28 104
rect 28 -104 44 104
rect -44 -123 44 -104
<< via2 >>
rect -28 -104 28 104
<< metal3 >>
rect -45 104 45 123
rect -45 -104 -28 104
rect 28 -104 45 104
rect -45 -123 45 -104
<< end >>
