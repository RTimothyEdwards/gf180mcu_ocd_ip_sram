magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< nwell >>
rect -174 -86 230 2202
<< pmos >>
rect 0 0 56 2116
<< pdiff >>
rect -88 2103 0 2116
rect -88 13 -75 2103
rect -29 13 0 2103
rect -88 0 0 13
rect 56 2103 144 2116
rect 56 13 85 2103
rect 131 13 144 2103
rect 56 0 144 13
<< pdiffc >>
rect -75 13 -29 2103
rect 85 13 131 2103
<< polysilicon >>
rect 0 2116 56 2160
rect 0 -44 56 0
<< metal1 >>
rect -75 2103 -29 2116
rect -75 0 -29 13
rect 85 2103 131 2116
rect 85 0 131 13
<< labels >>
flabel pdiffc -40 1058 -40 1058 0 FreeSans 186 0 0 0 S
flabel pdiffc 96 1058 96 1058 0 FreeSans 186 0 0 0 D
<< end >>
