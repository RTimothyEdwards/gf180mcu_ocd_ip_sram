magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< psubdiff >>
rect -62 81 62 95
rect -62 -81 -49 81
rect 49 -81 62 81
rect -62 -95 62 -81
<< psubdiffcont >>
rect -49 -81 49 81
<< metal1 >>
rect -56 81 56 89
rect -56 -81 -49 81
rect 49 -81 56 81
rect -56 -89 56 -81
<< end >>
