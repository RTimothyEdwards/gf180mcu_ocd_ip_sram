magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
use via1_x2_R270_3v256x8m81  via1_x2_R270_3v256x8m81_0
timestamp 1763766357
transform 1 0 0 0 1 0
box -8 0 75 215
use via2_x2_R270_3v256x8m81  via2_x2_R270_3v256x8m81_0
timestamp 1763766357
transform 1 0 0 0 1 0
box -9 0 75 215
<< end >>
