magic
tech gf180mcuD
magscale 1 10
timestamp 1763577663
<< metal1 >>
rect -45 1854 45 1874
rect -45 -1454 -26 1854
rect 26 -1454 45 1854
rect -45 -1474 45 -1454
<< via1 >>
rect -26 -1454 26 1854
<< metal2 >>
rect -45 1854 45 1874
rect -45 -1454 -26 1854
rect 26 -1454 45 1854
rect -45 -1474 45 -1454
<< end >>
