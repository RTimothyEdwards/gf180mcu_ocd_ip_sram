magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< nwell >>
rect -96 -86 96 86
<< nsubdiff >>
rect -72 23 72 46
rect -72 -23 -49 23
rect 49 -23 72 23
rect -72 -46 72 -23
<< nsubdiffcont >>
rect -49 -23 49 23
<< metal1 >>
rect -56 23 56 30
rect -56 -23 -49 23
rect 49 -23 56 23
rect -56 -30 56 -23
<< end >>
