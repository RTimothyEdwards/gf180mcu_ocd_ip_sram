magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal1 >>
rect -119 9844 119 9872
rect -119 -9844 -92 9844
rect 92 -9844 119 9844
rect -119 -9872 119 -9844
<< via1 >>
rect -92 -9844 92 9844
<< metal2 >>
rect -119 9844 119 9872
rect -119 -9844 -92 9844
rect 92 -9844 119 9844
rect -119 -9872 119 -9844
<< end >>
