magic
tech gf180mcuD
magscale 1 10
timestamp 1765917876
<< metal1 >>
rect 401 38753 447 38866
rect 401 37985 447 38098
rect 401 37541 447 37654
rect 401 36773 447 36886
rect 401 36329 447 36442
rect 401 35561 447 35674
rect 401 35117 447 35230
rect 401 34349 447 34462
rect 401 33905 447 34018
rect 401 33137 447 33250
rect 401 32693 447 32806
rect 401 31925 447 32038
rect 401 31481 447 31594
rect 401 30713 447 30826
rect 401 30269 447 30382
rect 401 29501 447 29614
rect 401 29057 447 29170
rect 401 28289 447 28402
rect 401 27845 447 27958
rect 401 27077 447 27190
rect 401 26633 447 26746
rect 401 25865 447 25978
rect 401 25421 447 25534
rect 401 24653 447 24766
rect 401 24209 447 24322
rect 401 23441 447 23554
rect 401 22997 447 23110
rect 401 22229 447 22342
rect 401 21785 447 21898
rect 401 21017 447 21130
rect 401 20573 447 20686
rect 401 19805 447 19918
rect 401 19361 447 19474
rect 401 18593 447 18706
rect 401 18149 447 18262
rect 401 17381 447 17494
rect 401 16937 447 17050
rect 401 16169 447 16282
rect 401 15725 447 15838
rect 401 14957 447 15070
rect 401 14513 447 14626
rect 401 13745 447 13858
rect 401 13301 447 13414
rect 401 12533 447 12646
rect 401 12089 447 12202
rect 401 11321 447 11434
rect 401 10877 447 10990
rect 401 10109 447 10222
rect 401 9665 447 9778
rect 401 8897 447 9010
rect 401 8453 447 8566
rect 401 7685 447 7798
rect 401 7241 447 7354
rect 401 6473 447 6586
rect 401 6029 447 6142
rect 401 5261 447 5374
rect 401 4817 447 4930
rect 401 4049 447 4162
rect 401 3605 447 3718
rect 401 2837 447 2950
rect 401 2393 447 2506
rect 401 1625 447 1738
rect 401 1181 447 1294
rect 401 413 447 526
<< metal2 >>
rect 734 129 854 229
rect 946 129 1066 229
rect 1170 129 1290 229
rect 1382 129 1502 229
rect 1606 129 1726 229
rect 1818 129 1938 229
rect 2042 129 2162 229
rect 2254 129 2374 229
rect 2478 129 2598 229
rect 2690 129 2810 229
rect 2914 129 3034 229
rect 3126 129 3246 229
rect 3350 129 3470 229
rect 3562 129 3682 229
rect 3786 129 3906 229
rect 3998 129 4118 229
rect 4642 129 4762 229
rect 4854 129 4974 229
rect 5078 129 5198 229
rect 5290 129 5410 229
rect 5514 129 5634 229
rect 5726 129 5846 229
rect 5950 129 6070 229
rect 6162 129 6282 229
rect 6386 129 6506 229
rect 6598 129 6718 229
rect 6822 129 6942 229
rect 7034 129 7154 229
rect 7258 129 7378 229
rect 7470 129 7590 229
rect 7694 129 7814 229
rect 7906 129 8026 229
rect 8550 129 8670 229
rect 8762 129 8882 229
rect 8986 129 9106 229
rect 9198 129 9318 229
rect 9422 129 9542 229
rect 9634 129 9754 229
rect 9858 129 9978 229
rect 10070 129 10190 229
rect 10294 129 10414 229
rect 10506 129 10626 229
rect 10730 129 10850 229
rect 10942 129 11062 229
rect 11166 129 11286 229
rect 11378 129 11498 229
rect 11602 129 11722 229
rect 11814 129 11934 229
rect 12458 129 12578 229
rect 12670 129 12790 229
rect 12894 129 13014 229
rect 13106 129 13226 229
rect 13330 129 13450 229
rect 13542 129 13662 229
rect 13766 129 13886 229
rect 13978 129 14098 229
rect 14202 129 14322 229
rect 14414 129 14534 229
rect 14638 129 14758 229
rect 14850 129 14970 229
rect 15074 129 15194 229
rect 15286 129 15406 229
rect 15510 129 15630 229
rect 15722 129 15842 229
use 018SRAM_cell1_2x_3v512x8m81  018SRAM_cell1_2x_3v512x8m81_0
array 0 7 -436 0 31 1212
timestamp 1764626446
transform -1 0 12924 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v512x8m81  018SRAM_cell1_2x_3v512x8m81_1
array 0 7 -436 0 31 1212
timestamp 1764626446
transform -1 0 5108 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v512x8m81  018SRAM_cell1_2x_3v512x8m81_2
array 0 7 436 0 31 1212
timestamp 1764626446
transform 1 0 600 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v512x8m81  018SRAM_cell1_2x_3v512x8m81_3
array 0 7 436 0 31 1212
timestamp 1764626446
transform 1 0 8416 0 1 0
box 30 103 570 1445
use 018SRAM_strap1_2x_3v512x8m81  018SRAM_strap1_2x_3v512x8m81_0
array 0 0 -420 0 31 1212
timestamp 1764693440
transform -1 0 12497 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_2x_3v512x8m81  018SRAM_strap1_2x_3v512x8m81_1
array 0 0 -420 0 31 1212
timestamp 1764693440
transform -1 0 773 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_2x_3v512x8m81  018SRAM_strap1_2x_3v512x8m81_2
array 0 0 -420 0 31 1212
timestamp 1764693440
transform -1 0 4681 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_2x_3v512x8m81  018SRAM_strap1_2x_3v512x8m81_3
array 0 0 -420 0 31 1212
timestamp 1764693440
transform -1 0 8589 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_2x_bndry_3v512x8m81  018SRAM_strap1_2x_bndry_3v512x8m81_0
array 0 0 420 0 31 1212
timestamp 1764625442
transform 1 0 15803 0 1 900
box 91 -797 511 545
<< labels >>
rlabel metal2 s 15780 170 15780 170 0 b[0]
rlabel metal2 s 15570 170 15570 170 0 bb[0]
rlabel metal2 s 15340 170 15340 170 0 bb[1]
rlabel metal2 s 15140 170 15140 170 0 b[1]
rlabel metal2 s 14910 170 14910 170 0 b[2]
rlabel metal2 s 14690 170 14690 170 0 bb[2]
rlabel metal2 s 14470 170 14470 170 0 bb[3]
rlabel metal2 s 14260 170 14260 170 0 b[3]
rlabel metal2 s 14030 170 14030 170 0 b[4]
rlabel metal2 s 13830 170 13830 170 0 bb[4]
rlabel metal2 s 13600 170 13600 170 0 bb[5]
rlabel metal2 s 13390 170 13390 170 0 b[5]
rlabel metal2 s 13160 170 13160 170 0 b[6]
rlabel metal2 s 12950 170 12950 170 0 bb[6]
rlabel metal2 s 12730 170 12730 170 0 bb[7]
rlabel metal2 s 12520 170 12520 170 0 b[7]
rlabel metal2 s 11870 170 11870 170 0 b[8]
rlabel metal2 s 11660 170 11660 170 0 bb[8]
rlabel metal2 s 11440 170 11440 170 0 bb[9]
rlabel metal2 s 11230 170 11230 170 0 b[9]
rlabel metal2 s 11000 170 11000 170 0 b[10]
rlabel metal2 s 10790 170 10790 170 0 bb[10]
rlabel metal2 s 10560 170 10560 170 0 bb[11]
rlabel metal2 s 10360 170 10360 170 0 b[11]
rlabel metal2 s 10130 170 10130 170 0 b[12]
rlabel metal2 s 9920 170 9920 170 0 bb[12]
rlabel metal2 s 9690 170 9690 170 0 bb[13]
rlabel metal2 s 9480 170 9480 170 0 b[13]
rlabel metal2 s 9260 170 9260 170 0 b[14]
rlabel metal2 s 9040 170 9040 170 0 bb[14]
rlabel metal2 s 8820 170 8820 170 0 bb[15]
rlabel metal2 s 8610 170 8610 170 0 b[15]
rlabel metal2 s 7960 170 7960 170 0 b[16]
rlabel metal2 s 7750 170 7750 170 0 bb[16]
rlabel metal2 s 7530 170 7530 170 0 bb[17]
rlabel metal2 s 7320 170 7320 170 0 b[17]
rlabel metal2 s 7090 170 7090 170 0 b[18]
rlabel metal2 s 6880 170 6880 170 0 bb[18]
rlabel metal2 s 6660 170 6660 170 0 bb[19]
rlabel metal2 s 6440 170 6440 170 0 b[19]
rlabel metal2 s 6220 170 6220 170 0 b[20]
rlabel metal2 s 6010 170 6010 170 0 bb[20]
rlabel metal2 s 5780 170 5780 170 0 bb[21]
rlabel metal2 s 5570 170 5570 170 0 b[21]
rlabel metal2 s 5350 170 5350 170 0 b[22]
rlabel metal2 s 5140 170 5140 170 0 bb[22]
rlabel metal2 s 4910 170 4910 170 0 bb[23]
rlabel metal2 s 4700 170 4700 170 0 b[23]
rlabel metal2 s 4060 170 4060 170 0 b[24]
rlabel metal2 s 3850 170 3850 170 0 bb[24]
rlabel metal2 s 3620 170 3620 170 0 bb[25]
rlabel metal2 s 3410 170 3410 170 0 b[25]
rlabel metal2 s 3180 170 3180 170 0 b[26]
rlabel metal2 s 2970 170 2970 170 0 bb[26]
rlabel metal2 s 2750 170 2750 170 0 bb[27]
rlabel metal2 s 2530 170 2530 170 0 b[27]
rlabel metal2 s 2310 170 2310 170 0 b[28]
rlabel metal2 s 2100 170 2100 170 0 bb[28]
rlabel metal2 s 1870 170 1870 170 0 bb[29]
rlabel metal2 s 1670 170 1670 170 0 b[29]
rlabel metal2 s 1440 170 1440 170 0 b[30]
rlabel metal2 s 1230 170 1230 170 0 bb[30]
rlabel metal2 s 1000 170 1000 170 0 bb[31]
rlabel metal2 s 790 170 790 170 0 b[31]
rlabel metal1 s 410 500 410 500 0 wl[0]
rlabel metal1 s 410 1260 410 1260 0 wl[1]
rlabel metal1 s 410 1720 410 1720 0 wl[2]
rlabel metal1 s 410 2930 410 2930 0 wl[4]
rlabel metal1 s 410 4130 410 4130 0 wl[6]
rlabel metal1 s 410 5350 410 5350 0 wl[8]
rlabel metal1 s 410 6550 410 6550 0 wl[10]
rlabel metal1 s 410 7760 410 7760 0 wl[12]
rlabel metal1 s 410 8530 410 8530 0 wl[13]
rlabel metal1 s 410 8980 410 8980 0 wl[14]
rlabel metal1 s 410 9750 410 9750 0 wl[15]
rlabel metal1 s 410 10190 410 10190 0 wl[16]
rlabel metal1 s 410 10950 410 10950 0 wl[17]
rlabel metal1 s 410 11400 410 11400 0 wl[18]
rlabel metal1 s 410 12170 410 12170 0 wl[19]
rlabel metal1 s 410 12620 410 12620 0 wl[20]
rlabel metal1 s 410 13380 410 13380 0 wl[21]
rlabel metal1 s 410 13830 410 13830 0 wl[22]
rlabel metal1 s 410 14590 410 14590 0 wl[23]
rlabel metal1 s 410 15040 410 15040 0 wl[24]
rlabel metal1 s 410 15810 410 15810 0 wl[25]
rlabel metal1 s 410 16250 410 16250 0 wl[26]
rlabel metal1 s 410 17020 410 17020 0 wl[27]
rlabel metal1 s 410 17470 410 17470 0 wl[28]
rlabel metal1 s 410 18230 410 18230 0 wl[29]
rlabel metal1 s 410 18670 410 18670 0 wl[30]
rlabel metal1 s 410 19440 410 19440 0 wl[31]
rlabel metal1 s 430 3660 430 3660 0 wl[5]
rlabel metal1 s 420 4890 420 4890 0 wl[7]
rlabel metal1 s 430 6090 430 6090 0 wl[9]
rlabel metal1 s 440 7310 440 7310 0 wl[11]
rlabel metal1 420 19860 420 19860 0 wl[32]
rlabel metal1 420 20620 420 20620 0 wl[33]
rlabel metal1 420 21070 420 21070 0 wl[34]
rlabel metal1 420 21850 420 21850 0 wl[35]
rlabel metal1 430 22280 430 22280 0 wl[36]
rlabel metal1 420 23050 420 23050 0 wl[37]
rlabel metal1 420 23500 420 23500 0 wl[38]
rlabel metal1 420 24260 420 24260 0 wl[39]
rlabel metal1 420 24710 420 24710 0 wl[40]
rlabel metal1 420 25470 420 25470 0 wl[41]
rlabel metal1 420 25920 420 25920 0 wl[42]
rlabel metal1 420 26690 420 26690 0 wl[43]
rlabel metal1 420 27130 420 27130 0 wl[44]
rlabel metal1 430 27900 430 27900 0 wl[45]
rlabel metal1 430 28340 430 28340 0 wl[46]
rlabel metal1 420 29110 420 29110 0 wl[47]
rlabel metal1 420 29560 420 29560 0 wl[48]
rlabel metal1 420 30320 420 30320 0 wl[49]
rlabel metal1 420 30770 420 30770 0 wl[50]
rlabel metal1 420 31540 420 31540 0 wl[51]
rlabel metal1 420 31980 420 31980 0 wl[52]
rlabel metal1 420 32750 420 32750 0 wl[53]
rlabel metal1 430 33190 430 33190 0 wl[54]
rlabel metal1 420 33960 420 33960 0 wl[55]
rlabel metal1 420 34410 420 34410 0 wl[56]
rlabel metal1 420 35170 420 35170 0 wl[57]
rlabel metal1 420 35620 420 35620 0 wl[58]
rlabel metal1 420 36380 420 36380 0 wl[59]
rlabel metal1 420 36830 420 36830 0 wl[60]
rlabel metal1 420 37590 420 37590 0 wl[61]
rlabel metal1 420 38040 420 38040 0 wl[62]
rlabel metal1 420 38810 420 38810 0 wl[63]
rlabel metal1 s 430 2450 430 2450 0 wl[3]
<< end >>
