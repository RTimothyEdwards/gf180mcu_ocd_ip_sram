magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal1 >>
rect -39 503 39 504
rect -44 502 42 503
rect -44 483 44 502
rect -44 -483 -26 483
rect 26 -483 44 483
rect -44 -503 44 -483
rect -35 -504 44 -503
<< via1 >>
rect -26 -483 26 483
<< metal2 >>
rect -44 483 44 502
rect -44 -483 -26 483
rect 26 -483 44 483
rect -44 -503 44 -483
<< end >>
