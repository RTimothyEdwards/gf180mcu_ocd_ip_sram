magic
tech gf180mcuD
magscale 1 10
timestamp 1765833452
<< polysilicon >>
rect 22200 20783 22260 20855
<< metal2 >>
rect 22231 172 22356 21009
<< metal3 >>
rect 5692 20808 22356 21008
rect 5727 173 22356 373
use 018SRAM_cell1_3v256x8m81  018SRAM_cell1_3v256x8m81_0
timestamp 1765833244
transform -1 0 22262 0 1 177
box 30 89 570 797
use 018SRAM_cell1_3v256x8m81  018SRAM_cell1_3v256x8m81_1
timestamp 1765833244
transform -1 0 22262 0 -1 21033
box 30 89 570 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_0
timestamp 1765833244
transform -1 0 16190 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_1
timestamp 1765833244
transform -1 0 15318 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_2
timestamp 1765833244
transform -1 0 15754 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_3
timestamp 1765833244
transform -1 0 14882 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_4
timestamp 1765833244
transform -1 0 18354 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_5
timestamp 1765833244
transform -1 0 18790 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_6
timestamp 1765833244
transform -1 0 19662 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_7
timestamp 1765833244
transform -1 0 19226 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_8
timestamp 1765833244
transform -1 0 20098 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_9
timestamp 1765833244
transform -1 0 20534 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_10
timestamp 1765833244
transform -1 0 20970 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_11
timestamp 1765833244
transform -1 0 21406 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_12
timestamp 1765833244
transform -1 0 17498 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_13
timestamp 1765833244
transform -1 0 17062 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_14
timestamp 1765833244
transform -1 0 16626 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_15
timestamp 1765833244
transform -1 0 6630 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_16
timestamp 1765833244
transform -1 0 10538 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_17
timestamp 1765833244
transform -1 0 10974 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_18
timestamp 1765833244
transform -1 0 11846 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_19
timestamp 1765833244
transform -1 0 11410 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_20
timestamp 1765833244
transform -1 0 12282 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_21
timestamp 1765833244
transform -1 0 12718 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_22
timestamp 1765833244
transform -1 0 13154 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_23
timestamp 1765833244
transform -1 0 13590 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_24
timestamp 1765833244
transform -1 0 9682 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_25
timestamp 1765833244
transform -1 0 9246 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_26
timestamp 1765833244
transform -1 0 8810 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_27
timestamp 1765833244
transform -1 0 8374 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_28
timestamp 1765833244
transform -1 0 7502 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_29
timestamp 1765833244
transform -1 0 7938 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_30
timestamp 1765833244
transform -1 0 7066 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_3v256x8m81  018SRAM_cell1_dummy_3v256x8m81_31
timestamp 1765833244
transform -1 0 14446 0 1 177
box 62 89 538 797
use 018SRAM_strap1_3v256x8m81  018SRAM_strap1_3v256x8m81_0
timestamp 1765833244
transform -1 0 17927 0 1 177
box 91 55 511 797
use 018SRAM_strap1_3v256x8m81  018SRAM_strap1_3v256x8m81_1
timestamp 1765833244
transform 1 0 21233 0 1 177
box 91 55 511 797
use 018SRAM_strap1_3v256x8m81  018SRAM_strap1_3v256x8m81_2
timestamp 1765833244
transform -1 0 14019 0 1 177
box 91 55 511 797
use 018SRAM_strap1_3v256x8m81  018SRAM_strap1_3v256x8m81_3
timestamp 1765833244
transform -1 0 10111 0 1 177
box 91 55 511 797
use 018SRAM_strap1_3v256x8m81  018SRAM_strap1_3v256x8m81_4
timestamp 1765833244
transform -1 0 6203 0 1 177
box 91 55 511 797
use 018SRAM_strap1_3v256x8m81  018SRAM_strap1_3v256x8m81_5
timestamp 1765833244
transform -1 0 6203 0 -1 21033
box 91 55 511 797
use array16_256_dummy_01_3v256x8m81  array16_256_dummy_01_3v256x8m81_0
timestamp 1764696963
transform 1 0 21594 0 1 673
box 98 171 638 20097
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_0
timestamp 1765833244
transform 1 0 22296 0 -1 17271
box -96 -124 67 124
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_1
timestamp 1765833244
transform 1 0 22296 0 -1 14847
box -96 -124 67 124
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_2
timestamp 1765833244
transform 1 0 22296 0 -1 11211
box -96 -124 67 124
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_3
timestamp 1765833244
transform 1 0 22296 0 -1 8787
box -96 -124 67 124
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_4
timestamp 1765833244
transform 1 0 22296 0 -1 6363
box -96 -124 67 124
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_5
timestamp 1765833244
transform 1 0 22296 0 -1 12423
box -96 -124 67 124
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_6
timestamp 1765833244
transform 1 0 22296 0 -1 9999
box -96 -124 67 124
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_7
timestamp 1765833244
transform 1 0 22296 0 -1 7575
box -96 -124 67 124
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_8
timestamp 1765833244
transform 1 0 22296 0 -1 5151
box -96 -124 67 124
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_9
timestamp 1765833244
transform 1 0 22296 0 -1 3939
box -96 -124 67 124
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_10
timestamp 1765833244
transform 1 0 22296 0 -1 1515
box -96 -124 67 124
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_11
timestamp 1765833244
transform 1 0 22296 0 -1 18483
box -96 -124 67 124
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_12
timestamp 1765833244
transform 1 0 22296 0 -1 16059
box -96 -124 67 124
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_13
timestamp 1765833244
transform 1 0 22296 0 -1 13635
box -96 -124 67 124
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_14
timestamp 1765833244
transform 1 0 22296 0 -1 2727
box -96 -124 67 124
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_15
timestamp 1765833244
transform 1 0 22296 0 -1 303
box -96 -124 67 124
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_16
timestamp 1765833244
transform 1 0 22296 0 -1 19695
box -96 -124 67 124
use M1_POLY24310591302019_3v256x8m81  M1_POLY24310591302019_3v256x8m81_0
timestamp 1765833244
transform 1 0 22295 0 1 20766
box -36 -80 36 78
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_0
timestamp 1765833244
transform 1 0 22294 0 -1 5153
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_1
timestamp 1765833244
transform 1 0 22294 0 -1 14849
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_2
timestamp 1765833244
transform 1 0 22294 0 -1 19693
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_3
timestamp 1765833244
transform 1 0 22294 0 -1 10001
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_4
timestamp 1765833244
transform 1 0 22294 0 -1 2727
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_5
timestamp 1765833244
transform 1 0 22294 0 -1 12425
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_6
timestamp 1765833244
transform 1 0 22294 0 -1 17273
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_7
timestamp 1765833244
transform 1 0 22294 0 -1 7577
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_8
timestamp 1765833244
transform 1 0 22294 0 -1 1513
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_9
timestamp 1765833244
transform 1 0 22294 0 -1 3937
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_10
timestamp 1765833244
transform 1 0 22294 0 -1 6361
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_11
timestamp 1765833244
transform 1 0 22294 0 -1 8785
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_12
timestamp 1765833244
transform 1 0 22294 0 -1 11209
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_13
timestamp 1765833244
transform 1 0 22294 0 -1 13633
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_14
timestamp 1765833244
transform 1 0 22294 0 -1 16057
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_15
timestamp 1765833244
transform 1 0 22294 0 -1 18481
box -43 -122 43 122
use M2_M1431059130208_3v256x8m81  M2_M1431059130208_3v256x8m81_0
timestamp 1765833244
transform 1 0 22294 0 1 297
box -34 -63 34 63
use M2_M14310591302018_3v256x8m81  M2_M14310591302018_3v256x8m81_0
timestamp 1765833244
transform 1 0 22295 0 1 20825
box -34 -99 34 99
use M3_M2431059130201_3v256x8m81  M3_M2431059130201_3v256x8m81_0
timestamp 1765833244
transform 1 0 22294 0 1 276
box -35 -63 35 63
use M3_M2431059130201_3v256x8m81  M3_M2431059130201_3v256x8m81_1
timestamp 1765833244
transform 1 0 22295 0 1 20937
box -35 -63 35 63
use new_dummyrow_unit_3v256x8m81  new_dummyrow_unit_3v256x8m81_0
timestamp 1765833452
transform 1 0 10971 0 -1 21210
box 2937 232 10773 974
use new_dummyrowunit01_3v256x8m81  new_dummyrowunit01_3v256x8m81_0
timestamp 1765833452
transform 1 0 3157 0 -1 21210
box 2935 232 10771 974
<< end >>
