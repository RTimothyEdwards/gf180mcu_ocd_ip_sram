magic
tech gf180mcuD
magscale 1 10
timestamp 1765833244
<< polysilicon >>
rect -123 23 123 48
rect -123 -23 -78 23
rect 78 -23 123 23
rect -123 -48 123 -23
<< polycontact >>
rect -78 -23 78 23
<< metal1 >>
rect -95 23 95 42
rect -95 -23 -78 23
rect 78 -23 95 23
rect -95 -42 95 -23
<< end >>
