magic
tech gf180mcuD
magscale 1 10
timestamp 1763580222
<< metal2 >>
rect -5 2486 151 4401
rect 346 2660 503 4904
rect 707 2486 864 4394
use M2_M14310591302097_512x8m81  M2_M14310591302097_512x8m81_0
timestamp 1763564386
transform 1 0 784 0 1 2869
box -70 -330 70 330
use M2_M14310591302097_512x8m81  M2_M14310591302097_512x8m81_1
timestamp 1763564386
transform 1 0 72 0 1 2869
box -70 -330 70 330
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_0
timestamp 1763564386
transform 1 0 424 0 1 4763
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_1
timestamp 1763564386
transform 1 0 786 0 1 3510
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_2
timestamp 1763564386
transform 1 0 786 0 1 4280
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_3
timestamp 1763564386
transform 1 0 74 0 1 4280
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_4
timestamp 1763564386
transform 1 0 74 0 1 3510
box -70 -113 70 113
use M3_M243105913020102_512x8m81  M3_M243105913020102_512x8m81_0
timestamp 1763564386
transform 1 0 424 0 1 2928
box -70 -243 70 243
<< end >>
