magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -1299 172 1299 198
rect -1299 -172 -1274 172
rect 1274 -172 1299 172
rect -1299 -198 1299 -172
<< via2 >>
rect -1274 -172 1274 172
<< metal3 >>
rect -1299 172 1299 198
rect -1299 -172 -1274 172
rect 1274 -172 1299 172
rect -1299 -198 1299 -172
<< end >>
