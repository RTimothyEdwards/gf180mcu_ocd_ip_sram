magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -330 440 330 447
rect -330 -540 -323 440
rect 323 -540 330 440
rect -330 -547 330 -540
<< via2 >>
rect -323 -540 323 440
<< metal3 >>
rect -330 440 330 447
rect -330 -540 -323 440
rect 323 -540 330 440
rect -330 -547 330 -540
<< end >>
