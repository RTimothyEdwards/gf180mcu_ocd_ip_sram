magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal1 >>
rect 2534 880 3234 910
rect 2534 519 3894 880
rect 2534 -140 3234 519
rect 3342 138 3599 170
rect 3342 58 3927 138
rect 3342 30 3597 58
<< metal3 >>
rect 2337 805 3047 945
rect 2337 595 21427 805
rect 2337 455 3047 595
rect 2337 -175 3531 315
use M2_M14310591302087_3v512x8m81  M2_M14310591302087_3v512x8m81_0
timestamp 1763765945
transform 1 0 2648 0 1 700
box -113 -243 113 243
use M2_M14310591302087_3v512x8m81  M2_M14310591302087_3v512x8m81_1
timestamp 1763765945
transform 1 0 3418 0 1 70
box -113 -243 113 243
use M3_M24310591302090_3v512x8m81  M3_M24310591302090_3v512x8m81_0
timestamp 1763765945
transform 1 0 3418 0 1 70
box -113 -243 113 243
use M3_M24310591302090_3v512x8m81  M3_M24310591302090_3v512x8m81_1
timestamp 1763765945
transform 1 0 2648 0 1 700
box -113 -243 113 243
<< properties >>
string path 25.225 0.500 16.695 0.500 
<< end >>
