magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -70 323 70 330
rect -70 -323 -63 323
rect 63 -323 70 323
rect -70 -330 70 -323
<< via2 >>
rect -63 -323 63 323
<< metal3 >>
rect -70 323 70 330
rect -70 -323 -63 323
rect 63 -323 70 323
rect -70 -330 70 -323
<< end >>
