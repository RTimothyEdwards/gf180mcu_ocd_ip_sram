magic
tech gf180mcuD
magscale 1 10
timestamp 1765833244
<< nwell >>
rect -596 -159 597 159
<< nsubdiff >>
rect -497 23 497 56
rect -497 -23 -466 23
rect 466 -23 497 23
rect -497 -56 497 -23
<< nsubdiffcont >>
rect -466 -23 466 23
<< metal1 >>
rect -483 23 483 42
rect -483 -23 -466 23
rect 466 -23 483 23
rect -483 -42 483 -23
<< end >>
