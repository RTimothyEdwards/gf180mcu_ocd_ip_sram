magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< psubdiff >>
rect -662 23 662 56
rect -662 -23 -632 23
rect 532 -23 662 23
rect -662 -56 662 -23
<< psubdiffcont >>
rect -632 -23 532 23
<< metal1 >>
rect -649 23 578 42
rect -649 -23 -632 23
rect 532 -23 578 23
rect -649 -42 578 -23
<< end >>
