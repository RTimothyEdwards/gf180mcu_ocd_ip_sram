magic
tech gf180mcuD
magscale 1 10
timestamp 1764700137
<< metal2 >>
rect 0 74 65 92
rect 0 17 3 74
rect 60 17 65 74
rect 0 0 65 17
<< via2 >>
rect 3 17 60 74
<< metal3 >>
rect 0 74 65 92
rect 0 17 3 74
rect 60 17 65 74
rect 0 0 65 17
<< end >>
