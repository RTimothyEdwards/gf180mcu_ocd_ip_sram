magic
tech gf180mcuD
magscale 1 10
timestamp 1764700137
<< error_p >>
rect -103 0 -57 112
rect 57 0 103 112
rect 217 0 263 112
<< nwell >>
rect -202 -86 362 198
<< pmos >>
rect -28 0 28 112
rect 132 0 188 112
<< pdiff >>
rect -116 98 -28 112
rect -116 13 -103 98
rect -57 13 -28 98
rect -116 0 -28 13
rect 28 98 132 112
rect 28 13 57 98
rect 103 13 132 98
rect 28 0 132 13
rect 188 98 276 112
rect 188 13 217 98
rect 263 13 276 98
rect 188 0 276 13
<< pdiffc >>
rect -103 13 -57 98
rect 57 13 103 98
rect 217 13 263 98
<< polysilicon >>
rect -28 112 28 156
rect 132 112 188 156
rect -28 -44 28 0
rect 132 -44 188 0
<< metal1 >>
rect -103 98 -57 112
rect -103 0 -57 13
rect 57 98 103 112
rect 57 0 103 13
rect 217 98 263 112
rect 217 0 263 13
<< labels >>
flabel pdiffc 80 56 80 56 0 FreeSans 186 0 0 0 D
flabel pdiffc -68 56 -68 56 0 FreeSans 186 0 0 0 S
flabel pdiffc 228 56 228 56 0 FreeSans 186 0 0 0 S
<< end >>
