magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< nwell >>
rect -174 -86 230 1952
<< pmos >>
rect 0 0 56 1866
<< pdiff >>
rect -88 1853 0 1866
rect -88 13 -75 1853
rect -29 13 0 1853
rect -88 0 0 13
rect 56 1853 144 1866
rect 56 13 85 1853
rect 131 13 144 1853
rect 56 0 144 13
<< pdiffc >>
rect -75 13 -29 1853
rect 85 13 131 1853
<< polysilicon >>
rect 0 1866 56 1910
rect 0 -44 56 0
<< metal1 >>
rect -75 1853 -29 1866
rect -75 0 -29 13
rect 85 1853 131 1866
rect 85 0 131 13
<< labels >>
flabel pdiffc -40 933 -40 933 0 FreeSans 186 0 0 0 S
flabel pdiffc 96 933 96 933 0 FreeSans 186 0 0 0 D
<< end >>
