magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect 1546 3580 3253 4708
rect 1521 3262 3287 3580
rect 1970 571 3163 644
<< psubdiff >>
rect 1395 4897 3523 5013
rect 3412 746 3523 4897
rect 1727 164 1838 291
rect 3412 242 3445 746
rect 3491 242 3523 746
rect 1727 163 1839 164
rect 3412 163 3523 242
rect 1727 48 3523 163
<< psubdiffcont >>
rect 3445 242 3491 746
<< polysilicon >>
rect 2217 4661 2594 4731
rect 2217 4546 2273 4661
rect 2377 4546 2433 4661
rect 2538 4546 2594 4661
rect 1734 3936 1790 4261
rect 1894 3936 1950 4261
rect 2380 3936 2436 4261
rect 2844 3936 2900 4261
rect 3004 3936 3060 4261
rect 1466 3605 1951 3644
rect 2844 3605 3303 3644
rect 1939 3259 2003 3318
rect 1784 3102 1873 3168
rect 1784 2765 1841 3102
rect 2107 3021 2164 3319
rect 2107 2986 2186 3021
rect 1946 2950 2186 2986
rect 1946 2940 2162 2950
rect 1946 2783 1999 2940
rect 1784 2674 1840 2765
rect 1944 2732 1999 2783
rect 2105 2767 2162 2940
rect 2271 2783 2324 3327
rect 2440 3325 2486 3327
rect 1944 2674 2000 2732
rect 2106 2674 2162 2767
rect 2266 2743 2324 2783
rect 2428 3176 2486 3325
rect 2428 3105 2530 3176
rect 2266 2674 2322 2743
rect 2428 2674 2484 3105
rect 2588 2986 2646 3327
rect 2750 3267 2884 3326
rect 2886 3098 2967 3168
rect 2588 2938 2806 2986
rect 2588 2674 2644 2938
rect 2749 2765 2806 2938
rect 2909 2769 2967 3098
rect 2750 2674 2806 2765
rect 2910 2674 2966 2769
rect 3071 2184 3127 2287
rect 1813 1712 1869 1716
rect 1973 1712 2029 1716
rect 2135 1712 2191 1716
rect 2295 1712 2351 1716
rect 2457 1712 2513 1716
rect 2617 1712 2673 1716
rect 2779 1712 2835 1716
rect 2939 1712 2995 1716
rect 1812 1704 2995 1712
rect 1812 1616 2993 1704
rect 2139 1121 2195 1259
rect 2120 1049 2355 1121
rect 2139 972 2195 1049
rect 2299 972 2355 1049
rect 2460 972 2516 1259
rect 2620 1238 2677 1259
rect 2781 1238 2837 1259
rect 2620 1197 2837 1238
rect 2620 1121 2676 1197
rect 2590 1049 2676 1121
rect 2941 1085 2997 1259
rect 2620 972 2676 1049
rect 2781 1040 2997 1085
rect 2781 972 2837 1040
rect 2941 972 2997 1040
<< metal1 >>
rect 1229 5555 1817 5623
rect 2153 5555 3150 5623
rect 1752 5476 1817 5555
rect 1752 5408 3150 5476
rect 1229 5234 3419 5331
rect 875 5085 3150 5153
rect 1291 4904 3517 5007
rect 2289 4776 2526 4829
rect 2370 4775 2437 4776
rect 1290 1465 1390 4718
rect 1670 4666 2317 4718
rect 1670 4292 1720 4666
rect 1979 4293 2025 4666
rect 2267 4298 2317 4666
rect 2371 4659 2437 4775
rect 2491 4666 3138 4718
rect 2491 4298 2541 4666
rect 2757 4298 2838 4666
rect 3087 4298 3138 4666
rect 1985 4292 2018 4293
rect 1664 4118 1726 4242
rect 1990 4118 2053 4242
rect 2294 4177 3141 4242
rect 1664 4053 2513 4118
rect 1664 3997 1726 4053
rect 1663 3712 1726 3997
rect 1444 1706 1495 3658
rect 1819 3636 1865 3747
rect 1985 3686 2033 4053
rect 2302 3636 2354 3769
rect 2767 3760 2814 4177
rect 1713 3584 2354 3636
rect 2465 3636 2517 3760
rect 2781 3759 2814 3760
rect 2927 3636 2979 3752
rect 3089 3713 3141 4177
rect 3095 3712 3127 3713
rect 2465 3584 3038 3636
rect 3250 3611 3441 3658
rect 1600 3516 1666 3517
rect 1584 3303 1666 3516
rect 1632 2901 1682 3023
rect 1713 2958 1764 3584
rect 2205 3516 2271 3517
rect 2536 3516 2601 3517
rect 1875 3264 1955 3482
rect 1632 2849 1757 2901
rect 1707 2633 1757 2849
rect 2029 2633 2082 3486
rect 2200 3303 2282 3516
rect 2158 3096 2327 3180
rect 2158 2941 2305 3028
rect 2375 2873 2425 3482
rect 2527 3303 2607 3516
rect 2477 3096 2630 3180
rect 2503 2941 2657 3028
rect 2350 2807 2425 2873
rect 2720 2808 2770 3481
rect 2827 3264 2908 3488
rect 2886 3105 2940 3172
rect 2987 2958 3038 3584
rect 3092 3516 3158 3517
rect 3092 3303 3173 3516
rect 3132 3025 3182 3173
rect 3131 2957 3182 3025
rect 3132 2901 3182 2957
rect 2350 2633 2400 2807
rect 2674 2754 2770 2808
rect 2996 2849 3182 2901
rect 2674 2633 2720 2754
rect 2996 2633 3042 2849
rect 1549 2187 1630 2633
rect 2029 2632 2054 2633
rect 1875 2271 1955 2387
rect 2200 2271 2282 2387
rect 2527 2271 2607 2387
rect 2834 2271 2881 2387
rect 1875 2206 2881 2271
rect 1892 1762 1972 2206
rect 2205 1762 2286 2206
rect 2519 1762 2599 2206
rect 2832 1762 2913 2206
rect 3178 2187 3259 2636
rect 3390 1706 3441 3611
rect 1444 1622 3441 1706
rect 1290 1362 1833 1465
rect 1733 157 1833 1362
rect 2224 1109 2270 1307
rect 2224 1061 2590 1109
rect 2047 381 2128 931
rect 2224 905 2270 1061
rect 2361 462 2441 931
rect 2046 378 2128 381
rect 2360 378 2441 462
rect 2674 378 2755 931
rect 2987 378 3068 931
rect 3418 746 3517 808
rect 3418 242 3445 746
rect 3491 242 3517 746
rect 3418 157 3517 242
rect 1733 54 3517 157
<< metal2 >>
rect 1754 5623 1816 5702
rect 2146 5623 2208 5734
rect 1702 5613 1816 5623
rect 1702 5555 1765 5613
rect 2135 5555 2208 5623
rect 1968 5408 2034 5476
rect 2659 5408 2722 5702
rect 3053 5623 3116 5747
rect 2795 5555 3116 5623
rect 1969 4718 2034 5408
rect 1968 4666 2034 4718
rect 2371 4659 2437 5153
rect 2795 4650 2860 5555
rect 1816 4242 1879 4524
rect 1449 4177 1879 4242
rect 1449 3173 1512 4177
rect 2293 4053 2359 4320
rect 2451 4053 2517 4320
rect 2926 4244 2991 4524
rect 2926 4176 3287 4244
rect 1449 3105 3122 3173
rect 1449 1616 1512 3105
rect 3221 3025 3287 4176
rect 1671 2957 3287 3025
rect 3221 1617 3287 2957
rect 1449 1551 1986 1616
rect 1924 1052 1986 1551
rect 2995 1549 3434 1617
rect 2370 1246 2435 1421
rect 2678 1246 2744 1421
rect 2992 1246 3058 1421
rect 2370 1178 2744 1246
rect 2842 1178 3058 1246
rect 2520 -137 2586 1178
rect 2842 -137 2907 1178
rect 3126 1052 3192 1549
<< metal3 >>
rect 1701 5555 2191 5623
rect 1701 5476 1766 5555
rect 1178 5408 1766 5476
rect -249 3068 3468 4974
rect -249 486 3504 2867
rect -249 -120 3504 381
use M1_NWELL06_512x8m81  M1_NWELL06_512x8m81_0
timestamp 1763476864
transform 1 0 2566 0 1 420
box -596 -159 597 159
use M1_NWELL_01_R90_512x8m81  M1_NWELL_01_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 1619 1 0 3421
box -159 -154 159 154
use M1_NWELL_01_R90_512x8m81  M1_NWELL_01_R90_512x8m81_1
timestamp 1763476864
transform 0 -1 3132 1 0 3421
box -159 -154 159 154
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_0
timestamp 1763476864
transform -1 0 2720 0 1 1664
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_1
timestamp 1763476864
transform -1 0 2925 0 1 1664
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_2
timestamp 1763476864
transform 1 0 3154 0 1 2232
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_3
timestamp 1763476864
transform -1 0 2092 0 1 1664
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_4
timestamp 1763476864
transform 1 0 1647 0 1 2231
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_5
timestamp 1763476864
transform 1 0 1880 0 1 1664
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_6
timestamp 1763476864
transform -1 0 2404 0 1 1664
box -67 -48 67 47
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1763476864
transform 1 0 2296 0 1 3138
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1763476864
transform 1 0 2181 0 1 2987
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_2
timestamp 1763476864
transform 1 0 1918 0 1 3288
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_3
timestamp 1763476864
transform 1 0 1495 0 1 3635
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_4
timestamp 1763476864
transform 1 0 1902 0 1 3138
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_5
timestamp 1763476864
transform 1 0 2633 0 1 2987
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_6
timestamp 1763476864
transform 1 0 2501 0 1 3138
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_7
timestamp 1763476864
transform 1 0 2906 0 1 3138
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_8
timestamp 1763476864
transform 1 0 2855 0 1 3290
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_9
timestamp 1763476864
transform 1 0 3273 0 1 3635
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_10
timestamp 1763476864
transform 1 0 2404 0 1 4701
box -36 -36 36 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_0
timestamp 1763476864
transform 1 0 2533 0 1 1085
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_1
timestamp 1763476864
transform 1 0 3052 0 1 1077
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_2
timestamp 1763476864
transform 1 0 2071 0 1 1085
box -62 -36 62 36
use M1_PSUB$$46555180_512x8m81  M1_PSUB$$46555180_512x8m81_0
timestamp 1763476864
transform 1 0 2407 0 1 4956
box -996 -58 996 57
use M1_PSUB$$46556204_512x8m81  M1_PSUB$$46556204_512x8m81_0
timestamp 1763476864
transform 1 0 1340 0 1 3185
box -56 -1829 56 1828
use M1_PSUB$$46557228_512x8m81  M1_PSUB$$46557228_512x8m81_0
timestamp 1763476864
transform 1 0 1561 0 1 1414
box -277 -58 277 58
use M1_PSUB$$46558252_512x8m81  M1_PSUB$$46558252_512x8m81_0
timestamp 1763476864
transform 1 0 2571 0 1 106
box -665 -58 665 57
use M1_PSUB_04_R90_512x8m81  M1_PSUB_04_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 1782 1 0 721
box -571 -56 571 55
use M3_M2$$43371564_512x8m81  M3_M2$$43371564_512x8m81_0
timestamp 1763476864
transform 1 0 3035 0 1 2224
box -119 -46 119 46
use M3_M2$$43371564_512x8m81  M3_M2$$43371564_512x8m81_1
timestamp 1763476864
transform 1 0 1769 0 1 2224
box -119 -46 119 46
use nmos_1p2$$45107244_512x8m81  nmos_1p2$$45107244_512x8m81_0
timestamp 1763476864
transform -1 0 2900 0 -1 1509
box -185 -44 527 255
use nmos_1p2$$46550060_512x8m81  nmos_1p2$$46550060_512x8m81_0
timestamp 1763476864
transform 1 0 2024 0 1 1757
box -299 -44 1060 309
use nmos_1p2$$46551084_512x8m81  nmos_1p2$$46551084_512x8m81_0
timestamp 1763476864
transform -1 0 2181 0 -1 1509
box -102 -44 130 255
use nmos_1p2$$46552108_512x8m81  nmos_1p2$$46552108_512x8m81_0
timestamp 1763476864
transform 1 0 1996 0 1 2321
box -301 -45 1060 363
use nmos_1p2$$46553132_512x8m81  nmos_1p2$$46553132_512x8m81_0
timestamp 1763476864
transform 1 0 3085 0 1 2321
box -102 -44 130 362
use nmos_1p2$$46553132_512x8m81  nmos_1p2$$46553132_512x8m81_1
timestamp 1763476864
transform 1 0 1638 0 1 2321
box -102 -44 130 362
use pmos_1p2$$46285868_512x8m81  pmos_1p2$$46285868_512x8m81_0
timestamp 1763476864
transform 1 0 2394 0 1 3686
box -188 -86 216 297
use pmos_1p2$$46286892_512x8m81  pmos_1p2$$46286892_512x8m81_0
timestamp 1763476864
transform 1 0 2287 0 1 4292
box -244 -86 481 297
use pmos_1p2$$46549036_512x8m81  pmos_1p2$$46549036_512x8m81_0
timestamp 1763476864
transform -1 0 2843 0 -1 931
box -328 -86 878 297
use pmos_1p2$$46896172_512x8m81  pmos_1p2$$46896172_512x8m81_0
timestamp 1763476864
transform 1 0 2206 0 1 3361
box -272 -86 613 170
use pmos_1p2$$46897196_512x8m81  pmos_1p2$$46897196_512x8m81_0
timestamp 1763476864
transform 1 0 1776 0 1 4292
box -216 -86 348 297
use pmos_1p2$$46897196_512x8m81  pmos_1p2$$46897196_512x8m81_1
timestamp 1763476864
transform 1 0 1776 0 1 3686
box -216 -86 348 297
use pmos_1p2$$46897196_512x8m81  pmos_1p2$$46897196_512x8m81_2
timestamp 1763476864
transform 1 0 2886 0 1 4292
box -216 -86 348 297
use pmos_1p2$$46897196_512x8m81  pmos_1p2$$46897196_512x8m81_3
timestamp 1763476864
transform 1 0 2886 0 1 3686
box -216 -86 348 297
use pmos_1p2$$46898220_512x8m81  pmos_1p2$$46898220_512x8m81_0
timestamp 1763476864
transform 1 0 1962 0 1 3361
box -188 -86 216 170
use pmos_1p2$$46898220_512x8m81  pmos_1p2$$46898220_512x8m81_1
timestamp 1763476864
transform 1 0 2763 0 1 3361
box -188 -86 216 170
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_0
timestamp 1763476864
transform 1 0 3436 0 1 578
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_1
timestamp 1763476864
transform 1 0 2683 0 1 1834
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_2
timestamp 1763476864
transform -1 0 2590 0 -1 1540
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_3
timestamp 1763476864
transform -1 0 2902 0 -1 1540
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_4
timestamp 1763476864
transform 1 0 2989 0 1 1834
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_5
timestamp 1763476864
transform 1 0 2370 0 1 1834
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_6
timestamp 1763476864
transform -1 0 2123 0 -1 1420
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_7
timestamp 1763476864
transform 1 0 1766 0 1 578
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_8
timestamp 1763476864
transform 1 0 1766 0 1 1141
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_9
timestamp 1763476864
transform 1 0 1750 0 1 1834
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_10
timestamp 1763476864
transform 1 0 2056 0 1 1834
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_11
timestamp 1763476864
transform 1 0 1890 0 1 3265
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_12
timestamp 1763476864
transform 1 0 2205 0 1 3305
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_13
timestamp 1763476864
transform 1 0 1592 0 1 3305
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_14
timestamp 1763476864
transform 1 0 2135 0 1 4357
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_15
timestamp 1763476864
transform 1 0 2536 0 1 3305
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_16
timestamp 1763476864
transform 1 0 2605 0 1 4357
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_17
timestamp 1763476864
transform 1 0 2828 0 1 3265
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_18
timestamp 1763476864
transform 1 0 3092 0 1 3305
box -9 0 73 215
use via1_2_x2_R90_512x8m81  via1_2_x2_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 2281 1 0 5555
box -9 0 73 215
use via1_2_x2_R270_512x8m81  via1_2_x2_R270_512x8m81_0
timestamp 1763476864
transform 0 1 2983 -1 0 380
box -9 0 75 215
use via1_2_x2_R270_512x8m81  via1_2_x2_R270_512x8m81_1
timestamp 1763476864
transform 0 1 1906 -1 0 380
box -9 0 75 215
use via1_2_x2_R270_512x8m81  via1_2_x2_R270_512x8m81_2
timestamp 1763476864
transform 0 1 2227 -1 0 380
box -9 0 75 215
use via1_512x8m81  via1_512x8m81_0
timestamp 1763476864
transform 1 0 2371 0 -1 4753
box 0 0 65 92
use via1_R90_512x8m81  via1_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 3154 1 0 2204
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_1
timestamp 1763476864
transform 0 -1 1740 1 0 2204
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_2
timestamp 1763476864
transform 0 -1 1764 1 0 2958
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_3
timestamp 1763476864
transform 0 -1 3077 1 0 3105
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_4
timestamp 1763476864
transform 0 -1 3197 1 0 2958
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_5
timestamp 1763476864
transform 0 -1 2516 1 0 4054
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_6
timestamp 1763476864
transform 0 1 2293 1 0 4174
box 0 0 65 89
use via1_R270_512x8m81  via1_R270_512x8m81_0
timestamp 1763476864
transform 0 -1 2047 -1 0 4733
box 0 0 67 89
use via1_R270_512x8m81  via1_R270_512x8m81_1
timestamp 1763476864
transform 0 1 2158 -1 0 3024
box 0 0 67 89
use via1_R270_512x8m81  via1_R270_512x8m81_2
timestamp 1763476864
transform 0 1 2235 -1 0 3172
box 0 0 67 89
use via1_R270_512x8m81  via1_R270_512x8m81_3
timestamp 1763476864
transform 0 -1 2450 -1 0 5152
box 0 0 67 89
use via1_R270_512x8m81  via1_R270_512x8m81_4
timestamp 1763476864
transform 0 -1 2842 -1 0 4718
box 0 0 67 89
use via1_R270_512x8m81  via1_R270_512x8m81_5
timestamp 1763476864
transform 0 1 2561 -1 0 3024
box 0 0 67 89
use via1_R270_512x8m81  via1_R270_512x8m81_6
timestamp 1763476864
transform 0 1 2359 -1 0 3024
box 0 0 67 89
use via1_R270_512x8m81  via1_R270_512x8m81_7
timestamp 1763476864
transform 0 1 2484 -1 0 3172
box 0 0 67 89
use via1_x2_512x8m81  via1_x2_512x8m81_0
timestamp 1763476864
transform -1 0 2907 0 1 712
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_1
timestamp 1763476864
transform 1 0 2993 0 1 1198
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_2
timestamp 1763476864
transform 1 0 2520 0 1 712
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_3
timestamp 1763476864
transform -1 0 2744 0 1 1198
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_4
timestamp 1763476864
transform -1 0 2434 0 1 1198
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_5
timestamp 1763476864
transform 1 0 1817 0 1 4302
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_6
timestamp 1763476864
transform 1 0 2926 0 1 4302
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_7
timestamp 1763476864
transform 1 0 2452 0 1 4302
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_8
timestamp 1763476864
transform -1 0 2358 0 1 4302
box -8 0 72 222
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 3191 1 0 1045
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_1
timestamp 1763476864
transform 0 -1 2139 1 0 1053
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_2
timestamp 1763476864
transform 0 -1 2110 1 0 5409
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_3
timestamp 1763476864
transform 0 -1 1843 1 0 5555
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_4
timestamp 1763476864
transform 0 -1 2713 1 0 5409
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_5
timestamp 1763476864
transform 0 -1 3147 1 0 5555
box -8 0 72 215
use via1_x2_R270_512x8m81  via1_x2_R270_512x8m81_0
timestamp 1763476864
transform 0 1 1878 -1 0 3172
box -8 0 75 215
use via1_x2_R270_512x8m81  via1_x2_R270_512x8m81_1
timestamp 1763476864
transform 0 1 2718 -1 0 3172
box -8 0 75 215
use via2_x2_R90_512x8m81  via2_x2_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 1394 1 0 5409
box -9 0 73 215
<< labels >>
rlabel metal3 s 825 3607 825 3607 4 vdd
port 1 nsew
rlabel metal3 s 872 1687 872 1687 4 vss
port 2 nsew
rlabel metal3 s 722 81 722 81 4 vdd
port 1 nsew
rlabel metal2 s 2553 -95 2553 -95 4 qp
port 3 nsew
rlabel metal2 s 2007 4921 2007 4921 4 d
port 5 nsew
rlabel metal2 s 2877 -95 2877 -95 4 qn
port 6 nsew
rlabel metal1 s 2416 5285 2416 5285 4 wep
port 7 nsew
rlabel metal1 s 2405 5597 2405 5597 4 db
port 4 nsew
rlabel metal1 s 3129 1682 3129 1682 4 se
port 8 nsew
rlabel metal1 s 1428 5106 1428 5106 4 pcb
port 9 nsew
rlabel metal1 s 2402 5446 2402 5446 4 d
port 5 nsew
rlabel metal2 s 2826 4921 2826 4921 4 db
port 4 nsew
<< end >>
