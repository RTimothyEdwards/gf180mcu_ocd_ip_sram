magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nwell >>
rect -722 -86 2732 1800
<< pmos >>
rect -548 0 -492 1714
rect -388 0 -332 1714
rect -227 0 -171 1714
rect -67 0 -11 1714
rect 94 0 150 1714
rect 254 0 310 1714
rect 415 0 471 1714
rect 575 0 631 1714
rect 736 0 792 1714
rect 896 0 952 1714
rect 1057 0 1113 1714
rect 1217 0 1273 1714
rect 1378 0 1434 1714
rect 1538 0 1594 1714
rect 1699 0 1755 1714
rect 1860 0 1916 1714
rect 2020 0 2076 1714
rect 2181 0 2237 1714
rect 2341 0 2397 1714
rect 2502 0 2558 1714
<< pdiff >>
rect -636 1701 -548 1714
rect -636 13 -623 1701
rect -577 13 -548 1701
rect -636 0 -548 13
rect -492 1701 -388 1714
rect -492 13 -463 1701
rect -417 13 -388 1701
rect -492 0 -388 13
rect -332 1701 -227 1714
rect -332 13 -303 1701
rect -257 13 -227 1701
rect -332 0 -227 13
rect -171 1701 -67 1714
rect -171 13 -142 1701
rect -96 13 -67 1701
rect -171 0 -67 13
rect -11 1701 94 1714
rect -11 13 18 1701
rect 64 13 94 1701
rect -11 0 94 13
rect 150 1701 254 1714
rect 150 13 179 1701
rect 225 13 254 1701
rect 150 0 254 13
rect 310 1701 415 1714
rect 310 13 339 1701
rect 385 13 415 1701
rect 310 0 415 13
rect 471 1701 575 1714
rect 471 13 500 1701
rect 546 13 575 1701
rect 471 0 575 13
rect 631 1701 736 1714
rect 631 13 660 1701
rect 706 13 736 1701
rect 631 0 736 13
rect 792 1701 896 1714
rect 792 13 821 1701
rect 867 13 896 1701
rect 792 0 896 13
rect 952 1701 1057 1714
rect 952 13 981 1701
rect 1027 13 1057 1701
rect 952 0 1057 13
rect 1113 1701 1217 1714
rect 1113 13 1142 1701
rect 1188 13 1217 1701
rect 1113 0 1217 13
rect 1273 1701 1378 1714
rect 1273 13 1302 1701
rect 1348 13 1378 1701
rect 1273 0 1378 13
rect 1434 1701 1538 1714
rect 1434 13 1463 1701
rect 1509 13 1538 1701
rect 1434 0 1538 13
rect 1594 1701 1699 1714
rect 1594 13 1623 1701
rect 1669 13 1699 1701
rect 1594 0 1699 13
rect 1755 1701 1860 1714
rect 1755 13 1784 1701
rect 1830 13 1860 1701
rect 1755 0 1860 13
rect 1916 1701 2020 1714
rect 1916 13 1945 1701
rect 1991 13 2020 1701
rect 1916 0 2020 13
rect 2076 1701 2181 1714
rect 2076 13 2105 1701
rect 2151 13 2181 1701
rect 2076 0 2181 13
rect 2237 1701 2341 1714
rect 2237 13 2266 1701
rect 2312 13 2341 1701
rect 2237 0 2341 13
rect 2397 1701 2502 1714
rect 2397 13 2426 1701
rect 2472 13 2502 1701
rect 2397 0 2502 13
rect 2558 1701 2646 1714
rect 2558 13 2587 1701
rect 2633 13 2646 1701
rect 2558 0 2646 13
<< pdiffc >>
rect -623 13 -577 1701
rect -463 13 -417 1701
rect -303 13 -257 1701
rect -142 13 -96 1701
rect 18 13 64 1701
rect 179 13 225 1701
rect 339 13 385 1701
rect 500 13 546 1701
rect 660 13 706 1701
rect 821 13 867 1701
rect 981 13 1027 1701
rect 1142 13 1188 1701
rect 1302 13 1348 1701
rect 1463 13 1509 1701
rect 1623 13 1669 1701
rect 1784 13 1830 1701
rect 1945 13 1991 1701
rect 2105 13 2151 1701
rect 2266 13 2312 1701
rect 2426 13 2472 1701
rect 2587 13 2633 1701
<< polysilicon >>
rect -548 1714 -492 1758
rect -388 1714 -332 1758
rect -227 1714 -171 1758
rect -67 1714 -11 1758
rect 94 1714 150 1758
rect 254 1714 310 1758
rect 415 1714 471 1758
rect 575 1714 631 1758
rect 736 1714 792 1758
rect 896 1714 952 1758
rect 1057 1714 1113 1758
rect 1217 1714 1273 1758
rect 1378 1714 1434 1758
rect 1538 1714 1594 1758
rect 1699 1714 1755 1758
rect 1860 1714 1916 1758
rect 2020 1714 2076 1758
rect 2181 1714 2237 1758
rect 2341 1714 2397 1758
rect 2502 1714 2558 1758
rect -548 -44 -492 0
rect -388 -44 -332 0
rect -227 -44 -171 0
rect -67 -44 -11 0
rect 94 -44 150 0
rect 254 -44 310 0
rect 415 -44 471 0
rect 575 -44 631 0
rect 736 -44 792 0
rect 896 -44 952 0
rect 1057 -44 1113 0
rect 1217 -44 1273 0
rect 1378 -44 1434 0
rect 1538 -44 1594 0
rect 1699 -44 1755 0
rect 1860 -44 1916 0
rect 2020 -44 2076 0
rect 2181 -44 2237 0
rect 2341 -44 2397 0
rect 2502 -44 2558 0
<< metal1 >>
rect -623 1701 -577 1714
rect -623 0 -577 13
rect -463 1701 -417 1714
rect -463 0 -417 13
rect -303 1701 -257 1714
rect -303 0 -257 13
rect -142 1701 -96 1714
rect -142 0 -96 13
rect 18 1701 64 1714
rect 18 0 64 13
rect 179 1701 225 1714
rect 179 0 225 13
rect 339 1701 385 1714
rect 339 0 385 13
rect 500 1701 546 1714
rect 500 0 546 13
rect 660 1701 706 1714
rect 660 0 706 13
rect 821 1701 867 1714
rect 821 0 867 13
rect 981 1701 1027 1714
rect 981 0 1027 13
rect 1142 1701 1188 1714
rect 1142 0 1188 13
rect 1302 1701 1348 1714
rect 1302 0 1348 13
rect 1463 1701 1509 1714
rect 1463 0 1509 13
rect 1623 1701 1669 1714
rect 1623 0 1669 13
rect 1784 1701 1830 1714
rect 1784 0 1830 13
rect 1945 1701 1991 1714
rect 1945 0 1991 13
rect 2105 1701 2151 1714
rect 2105 0 2151 13
rect 2266 1701 2312 1714
rect 2266 0 2312 13
rect 2426 1701 2472 1714
rect 2426 0 2472 13
rect 2587 1701 2633 1714
rect 2587 0 2633 13
<< labels >>
flabel pdiffc 1005 857 1005 857 0 FreeSans 186 0 0 0 S
flabel pdiffc 856 857 856 857 0 FreeSans 186 0 0 0 D
flabel pdiffc 696 857 696 857 0 FreeSans 186 0 0 0 S
flabel pdiffc 535 857 535 857 0 FreeSans 186 0 0 0 D
flabel pdiffc 374 857 374 857 0 FreeSans 186 0 0 0 S
flabel pdiffc 214 857 214 857 0 FreeSans 186 0 0 0 D
flabel pdiffc 53 857 53 857 0 FreeSans 186 0 0 0 S
flabel pdiffc -107 857 -107 857 0 FreeSans 186 0 0 0 D
flabel pdiffc -268 857 -268 857 0 FreeSans 186 0 0 0 S
flabel pdiffc -428 857 -428 857 0 FreeSans 186 0 0 0 D
flabel pdiffc -588 857 -588 857 0 FreeSans 186 0 0 0 S
flabel pdiffc 1153 857 1153 857 0 FreeSans 186 0 0 0 D
flabel pdiffc 1314 857 1314 857 0 FreeSans 186 0 0 0 S
flabel pdiffc 1474 857 1474 857 0 FreeSans 186 0 0 0 D
flabel pdiffc 1635 857 1635 857 0 FreeSans 186 0 0 0 S
flabel pdiffc 1795 857 1795 857 0 FreeSans 186 0 0 0 D
flabel pdiffc 1956 857 1956 857 0 FreeSans 186 0 0 0 S
flabel pdiffc 2116 857 2116 857 0 FreeSans 186 0 0 0 D
flabel pdiffc 2277 857 2277 857 0 FreeSans 186 0 0 0 S
flabel pdiffc 2598 857 2598 857 0 FreeSans 186 0 0 0 S
flabel pdiffc 2436 857 2436 857 0 FreeSans 186 0 0 0 D
<< end >>
