magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal1 >>
rect -1299 170 1299 198
rect -1299 -170 -1272 170
rect 1272 -170 1299 170
rect -1299 -198 1299 -170
<< via1 >>
rect -1272 -170 1272 170
<< metal2 >>
rect -1299 170 1299 198
rect -1299 -170 -1272 170
rect 1272 -170 1299 170
rect -1299 -198 1299 -170
<< end >>
