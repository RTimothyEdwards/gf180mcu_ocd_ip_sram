magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< error_s >>
rect 341 1390 371 1510
rect 340 1166 371 1390
rect 340 557 371 571
<< nwell >>
rect 341 1390 1141 1714
rect 2 557 251 1390
rect 340 557 1141 1390
<< psubdiff >>
rect 77 362 170 396
rect 77 202 100 362
rect 146 202 170 362
rect 77 167 170 202
<< nsubdiff >>
rect 77 1267 170 1292
rect 77 816 100 1267
rect 146 816 170 1267
rect 77 710 170 816
<< psubdiffcont >>
rect 100 202 146 362
<< nsubdiffcont >>
rect 100 816 146 1267
<< polysilicon >>
rect 527 1637 583 1813
rect 886 1768 942 1814
rect 886 1722 1166 1768
rect 527 1439 583 1488
rect 262 1397 583 1439
rect 887 1415 941 1484
rect 887 1360 963 1415
rect 1107 1233 1166 1722
rect 886 1185 1166 1233
rect 886 1077 942 1185
rect 372 604 428 618
rect 532 604 588 618
rect 372 508 716 604
rect 886 520 1110 562
rect 372 415 428 508
rect 532 415 588 508
rect 886 395 942 520
<< metal1 >>
rect 442 2004 1030 2077
rect 442 1481 523 2004
rect 251 1426 336 1427
rect 251 1362 523 1426
rect 83 1267 366 1285
rect 83 816 100 1267
rect 146 816 366 1267
rect 83 662 366 816
rect 82 362 366 454
rect 82 208 100 362
rect 83 202 100 208
rect 146 212 366 362
rect 442 247 523 1362
rect 599 1341 680 1615
rect 598 1227 680 1341
rect 802 598 883 1947
rect 959 1481 1030 2004
rect 1098 1681 1179 1765
rect 938 1348 1150 1431
rect 1094 1284 1150 1348
rect 1094 1200 1183 1284
rect 609 515 883 598
rect 801 514 883 515
rect 146 202 163 212
rect 83 173 163 202
rect 802 138 883 514
rect 938 331 1015 1143
rect 1094 526 1150 1200
rect 938 247 1032 331
rect 938 148 1015 247
<< metal3 >>
rect 0 1563 1184 2041
rect 0 754 1184 1390
rect -63 0 1184 634
use M1_POLY2_155_512x8m81  M1_POLY2_155_512x8m81_0
timestamp 1763476864
transform 1 0 648 0 1 557
box -67 -48 67 47
use M1_POLY2_155_512x8m81  M1_POLY2_155_512x8m81_1
timestamp 1763476864
transform 1 0 1110 0 1 568
box -67 -48 67 47
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_0
timestamp 1763476864
transform 1 0 1136 0 1 1707
box -36 -126 60 122
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1763476864
transform 1 0 977 0 1 1390
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1763476864
transform 1 0 291 0 1 1447
box -36 -36 36 36
use M1_PSUB$$45110316_512x8m81  M1_PSUB$$45110316_512x8m81_0
timestamp 1763476864
transform 1 0 214 0 1 1926
box -110 -58 111 57
use M2_M1$$43379756_153_512x8m81  M2_M1$$43379756_153_512x8m81_0
timestamp 1763476864
transform 1 0 639 0 1 1066
box -44 -275 44 275
use M2_M1$$43380780_152_512x8m81  M2_M1$$43380780_152_512x8m81_0
timestamp 1763476864
transform 1 0 127 0 1 1069
box -44 -198 45 198
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_0
timestamp 1763476864
transform 1 0 1139 0 1 1696
box -44 -123 44 122
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_1
timestamp 1763476864
transform 1 0 1138 0 1 1309
box -44 -123 44 122
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_2
timestamp 1763476864
transform 1 0 994 0 1 271
box -44 -123 44 122
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_3
timestamp 1763476864
transform 1 0 124 0 1 331
box -44 -123 44 122
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_4
timestamp 1763476864
transform 1 0 639 0 1 1817
box -44 -123 44 122
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_5
timestamp 1763476864
transform 1 0 123 0 1 1817
box -44 -123 44 122
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_6
timestamp 1763476864
transform 1 0 639 0 1 331
box -44 -123 44 122
use M3_M2$$43368492_151_512x8m81  M3_M2$$43368492_151_512x8m81_0
timestamp 1763476864
transform 1 0 639 0 1 331
box -45 -123 45 123
use M3_M2$$43368492_151_512x8m81  M3_M2$$43368492_151_512x8m81_1
timestamp 1763476864
transform 1 0 124 0 1 331
box -45 -123 45 123
use M3_M2$$47108140_149_512x8m81  M3_M2$$47108140_149_512x8m81_0
timestamp 1763476864
transform 1 0 127 0 1 1069
box -45 -198 45 198
use M3_M2$$47108140_149_512x8m81  M3_M2$$47108140_149_512x8m81_1
timestamp 1763476864
transform 1 0 123 0 1 1817
box -45 -198 45 198
use M3_M2$$47108140_149_512x8m81  M3_M2$$47108140_149_512x8m81_2
timestamp 1763476864
transform 1 0 639 0 1 1817
box -45 -198 45 198
use M3_M2$$47333420_150_512x8m81  M3_M2$$47333420_150_512x8m81_0
timestamp 1763476864
transform 1 0 639 0 1 1066
box -45 -275 45 275
use nmos_1p2$$47329324_512x8m81  nmos_1p2$$47329324_512x8m81_0
timestamp 1763476864
transform 1 0 414 0 1 206
box -130 -44 262 213
use nmos_1p2_157_512x8m81  nmos_1p2_157_512x8m81_0
timestamp 1763476864
transform 1 0 900 0 1 142
box -102 -44 130 255
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_0
timestamp 1763476864
transform 1 0 527 0 -1 1945
box -88 -44 144 133
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_1
timestamp 1763476864
transform 1 0 886 0 -1 1945
box -88 -44 144 133
use pmos_1p2$$47331372_512x8m81  pmos_1p2$$47331372_512x8m81_0
timestamp 1763476864
transform 1 0 414 0 1 657
box -216 -86 348 509
use pmos_1p2_160_512x8m81  pmos_1p2_160_512x8m81_0
timestamp 1763476864
transform 1 0 900 0 1 825
box -188 -86 216 297
use pmos_1p2_161_512x8m81  pmos_1p2_161_512x8m81_0
timestamp 1763476864
transform 1 0 900 0 -1 1615
box -188 -86 216 175
use pmos_1p2_161_512x8m81  pmos_1p2_161_512x8m81_1
timestamp 1763476864
transform 1 0 541 0 -1 1615
box -188 -86 216 175
<< labels >>
rlabel metal3 s 141 1808 141 1808 4 vss
port 1 nsew
rlabel metal3 s 92 256 92 256 4 vss
port 1 nsew
rlabel metal3 s 109 1048 109 1048 4 vdd
port 2 nsew
rlabel metal1 s 1138 1723 1138 1723 4 enb
port 3 nsew
rlabel metal1 s 483 289 483 289 4 ab
port 5 nsew
rlabel metal1 s 991 289 991 289 4 a
port 6 nsew
rlabel metal1 s 1142 1242 1142 1242 4 en
port 4 nsew
<< end >>
