magic
tech gf180mcuD
magscale 1 10
timestamp 1764700137
<< psubdiff >>
rect -627 23 594 54
rect -627 -23 -594 23
rect 561 -23 594 23
rect -627 -54 594 -23
<< psubdiffcont >>
rect -594 -23 561 23
<< metal1 >>
rect -613 23 613 40
rect -613 -23 -594 23
rect 561 -23 613 23
rect -613 -40 613 -23
<< end >>
