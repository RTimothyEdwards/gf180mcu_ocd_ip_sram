magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal1 >>
rect -107 26 107 46
rect -107 -26 -89 26
rect 89 -26 107 26
rect -107 -46 107 -26
<< via1 >>
rect -89 -26 89 26
<< metal2 >>
rect -107 26 107 46
rect -107 -26 -89 26
rect 89 -26 107 26
rect -107 -46 107 -26
<< end >>
