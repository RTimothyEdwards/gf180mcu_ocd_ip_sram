magic
tech gf180mcuD
magscale 1 10
timestamp 1763482574
<< error_s >>
rect 9113 20520 9123 20523
rect 9159 20520 9169 20523
rect 9358 20520 9368 20523
rect 9404 20520 9414 20523
rect 50173 20520 50183 20523
rect 50219 20520 50229 20523
rect 50418 20520 50428 20523
rect 50464 20520 50474 20523
rect 58234 20516 58244 20519
rect 58280 20516 58290 20519
rect 57987 20512 57997 20515
rect 58033 20512 58043 20515
rect 16877 20506 16887 20509
rect 16923 20506 16933 20509
rect 17125 20506 17135 20509
rect 17171 20506 17181 20509
rect 9113 20073 9123 20076
rect 9159 20073 9169 20076
rect 9358 20073 9368 20076
rect 9404 20073 9414 20076
rect 50173 20073 50183 20076
rect 50219 20073 50229 20076
rect 50418 20073 50428 20076
rect 50464 20073 50474 20076
rect 58234 20069 58244 20072
rect 58280 20069 58290 20072
rect 57987 20065 57997 20068
rect 58033 20065 58043 20068
rect 16877 20059 16887 20062
rect 16923 20059 16933 20062
rect 17125 20059 17135 20062
rect 17171 20059 17181 20062
rect 9113 19768 9123 19771
rect 9159 19768 9169 19771
rect 9358 19768 9368 19771
rect 9404 19768 9414 19771
rect 50173 19768 50183 19771
rect 50219 19768 50229 19771
rect 50418 19768 50428 19771
rect 50464 19768 50474 19771
rect 58234 19764 58244 19767
rect 58280 19764 58290 19767
rect 57987 19760 57997 19763
rect 58033 19760 58043 19763
rect 16877 19754 16887 19757
rect 16923 19754 16933 19757
rect 17125 19754 17135 19757
rect 17171 19754 17181 19757
rect 9113 19163 9123 19166
rect 9159 19163 9169 19166
rect 9358 19163 9368 19166
rect 9404 19163 9414 19166
rect 50173 19163 50183 19166
rect 50219 19163 50229 19166
rect 50418 19163 50428 19166
rect 50464 19163 50474 19166
rect 58234 19159 58244 19162
rect 58280 19159 58290 19162
rect 57987 19155 57997 19158
rect 58033 19155 58043 19158
rect 16877 19149 16887 19152
rect 16923 19149 16933 19152
rect 17125 19149 17135 19152
rect 17171 19149 17181 19152
<< metal1 >>
rect 1620 23625 1690 24201
rect 16965 23631 17035 24207
rect 42674 23618 42820 24194
rect 50470 23787 50617 24210
rect 58031 23620 58101 24193
<< metal2 >>
rect 5532 24523 5602 24645
rect 13342 24583 13412 24655
rect 5415 24453 5602 24523
rect 13197 24513 13412 24583
rect 46613 24523 46683 24803
rect 54433 24523 54503 24738
rect 5415 24088 5485 24453
rect 13197 24091 13267 24513
rect 46528 24453 46683 24523
rect 54388 24453 54503 24523
rect 1338 19148 1408 22814
rect 9151 22643 9221 23101
rect 9151 22573 9418 22643
rect 9353 22340 9418 22573
rect 17248 22359 17318 23028
rect 17119 22289 17318 22359
rect 42407 19165 42477 24332
rect 46528 24096 46598 24453
rect 50221 22656 50291 24330
rect 54388 24089 54458 24453
rect 50221 22586 50479 22656
rect 50414 22322 50479 22586
rect 58313 22375 58383 22814
rect 58231 22305 58383 22375
<< metal3 >>
rect 32887 10510 33562 11748
rect 19282 10453 33562 10510
rect 19282 10152 33378 10453
rect 29045 10143 33378 10152
rect 29045 9610 32183 10143
rect 28805 4614 35862 5174
use M2_M14310591302025_512x8m81  M2_M14310591302025_512x8m81_0
timestamp 1763476864
transform 0 1 13153 -1 0 24111
box -34 -85 34 135
use M2_M14310591302025_512x8m81  M2_M14310591302025_512x8m81_1
timestamp 1763476864
transform 0 1 46496 -1 0 24100
box -34 -85 34 135
use M2_M14310591302025_512x8m81  M2_M14310591302025_512x8m81_2
timestamp 1763476864
transform 0 1 54317 -1 0 24124
box -34 -85 34 135
use M2_M14310591302025_512x8m81  M2_M14310591302025_512x8m81_3
timestamp 1763476864
transform 0 1 5426 -1 0 24122
box -34 -85 34 135
use M2_M14310591302076_512x8m81  M2_M14310591302076_512x8m81_0
timestamp 1763476864
transform -1 0 50558 0 1 23926
box -34 -281 34 281
use M2_M14310591302076_512x8m81  M2_M14310591302076_512x8m81_1
timestamp 1763476864
transform -1 0 58066 0 1 23906
box -34 -281 34 281
use M2_M14310591302076_512x8m81  M2_M14310591302076_512x8m81_2
timestamp 1763476864
transform -1 0 42748 0 1 23916
box -34 -281 34 281
use M2_M14310591302076_512x8m81  M2_M14310591302076_512x8m81_3
timestamp 1763476864
transform 1 0 9458 0 1 23928
box -34 -281 34 281
use M2_M14310591302076_512x8m81  M2_M14310591302076_512x8m81_4
timestamp 1763476864
transform 1 0 1655 0 1 23926
box -34 -281 34 281
use M2_M14310591302076_512x8m81  M2_M14310591302076_512x8m81_5
timestamp 1763476864
transform 1 0 17002 0 1 23916
box -34 -281 34 281
use M3_M24310591302077_512x8m81  M3_M24310591302077_512x8m81_0
timestamp 1763476864
transform 1 0 9141 0 1 19467
box -35 -304 35 304
use M3_M24310591302077_512x8m81  M3_M24310591302077_512x8m81_1
timestamp 1763476864
transform 1 0 17153 0 1 19453
box -35 -304 35 304
use M3_M24310591302077_512x8m81  M3_M24310591302077_512x8m81_2
timestamp 1763476864
transform 1 0 16905 0 1 19453
box -35 -304 35 304
use M3_M24310591302077_512x8m81  M3_M24310591302077_512x8m81_3
timestamp 1763476864
transform 1 0 50446 0 1 19467
box -35 -304 35 304
use M3_M24310591302077_512x8m81  M3_M24310591302077_512x8m81_4
timestamp 1763476864
transform 1 0 50201 0 1 19467
box -35 -304 35 304
use M3_M24310591302077_512x8m81  M3_M24310591302077_512x8m81_5
timestamp 1763476864
transform 1 0 58262 0 1 19463
box -35 -304 35 304
use M3_M24310591302077_512x8m81  M3_M24310591302077_512x8m81_6
timestamp 1763476864
transform 1 0 58015 0 1 19459
box -35 -304 35 304
use M3_M24310591302077_512x8m81  M3_M24310591302077_512x8m81_7
timestamp 1763476864
transform 1 0 9386 0 1 19467
box -35 -304 35 304
use M3_M24310591302078_512x8m81  M3_M24310591302078_512x8m81_0
timestamp 1763476864
transform 1 0 9141 0 1 20298
box -35 -225 35 225
use M3_M24310591302078_512x8m81  M3_M24310591302078_512x8m81_1
timestamp 1763476864
transform 1 0 17153 0 1 20284
box -35 -225 35 225
use M3_M24310591302078_512x8m81  M3_M24310591302078_512x8m81_2
timestamp 1763476864
transform 1 0 16905 0 1 20284
box -35 -225 35 225
use M3_M24310591302078_512x8m81  M3_M24310591302078_512x8m81_3
timestamp 1763476864
transform 1 0 50446 0 1 20298
box -35 -225 35 225
use M3_M24310591302078_512x8m81  M3_M24310591302078_512x8m81_4
timestamp 1763476864
transform 1 0 50201 0 1 20298
box -35 -225 35 225
use M3_M24310591302078_512x8m81  M3_M24310591302078_512x8m81_5
timestamp 1763476864
transform 1 0 58262 0 1 20294
box -35 -225 35 225
use M3_M24310591302078_512x8m81  M3_M24310591302078_512x8m81_6
timestamp 1763476864
transform 1 0 58015 0 1 20290
box -35 -225 35 225
use M3_M24310591302078_512x8m81  M3_M24310591302078_512x8m81_7
timestamp 1763476864
transform 1 0 9386 0 1 20298
box -35 -225 35 225
use M3_M24310591302079_512x8m81  M3_M24310591302079_512x8m81_0
timestamp 1763476864
transform 1 0 42441 0 1 19832
box -35 -635 35 635
use M3_M24310591302079_512x8m81  M3_M24310591302079_512x8m81_1
timestamp 1763476864
transform 1 0 1373 0 1 19852
box -35 -635 35 635
<< properties >>
string path 205.755 34.960 256.160 34.960 
<< end >>
