magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< error_s >>
rect 16877 20656 16887 20659
rect 16923 20656 16933 20659
rect 17125 20656 17135 20659
rect 17171 20656 17181 20659
rect 9113 20650 9123 20653
rect 9159 20650 9169 20653
rect 9358 20650 9368 20653
rect 9404 20650 9414 20653
rect 50174 20647 50184 20650
rect 50220 20647 50230 20650
rect 50419 20647 50429 20650
rect 50465 20647 50475 20650
rect 58234 20646 58244 20649
rect 58280 20646 58290 20649
rect 57987 20642 57997 20645
rect 58033 20642 58043 20645
rect 16877 20209 16887 20212
rect 16923 20209 16933 20212
rect 17125 20209 17135 20212
rect 17171 20209 17181 20212
rect 9113 20203 9123 20206
rect 9159 20203 9169 20206
rect 9358 20203 9368 20206
rect 9404 20203 9414 20206
rect 50174 20200 50184 20203
rect 50220 20200 50230 20203
rect 50419 20200 50429 20203
rect 50465 20200 50475 20203
rect 58234 20199 58244 20202
rect 58280 20199 58290 20202
rect 57987 20195 57997 20198
rect 58033 20195 58043 20198
rect 16877 19904 16887 19907
rect 16923 19904 16933 19907
rect 17125 19904 17135 19907
rect 17171 19904 17181 19907
rect 9113 19898 9123 19901
rect 9159 19898 9169 19901
rect 9358 19898 9368 19901
rect 9404 19898 9414 19901
rect 50174 19895 50184 19898
rect 50220 19895 50230 19898
rect 50419 19895 50429 19898
rect 50465 19895 50475 19898
rect 58234 19894 58244 19897
rect 58280 19894 58290 19897
rect 57987 19890 57997 19893
rect 58033 19890 58043 19893
rect 16877 19299 16887 19302
rect 16923 19299 16933 19302
rect 17125 19299 17135 19302
rect 17171 19299 17181 19302
rect 9113 19293 9123 19296
rect 9159 19293 9169 19296
rect 9358 19293 9368 19296
rect 9404 19293 9414 19296
rect 50174 19290 50184 19293
rect 50220 19290 50230 19293
rect 50419 19290 50429 19293
rect 50465 19290 50475 19293
rect 58234 19289 58244 19292
rect 58280 19289 58290 19292
rect 57987 19285 57997 19288
rect 58033 19285 58043 19288
<< metal1 >>
rect 1620 23625 1690 24201
rect 16965 23631 17035 24207
rect 42674 23618 42820 24194
rect 50470 23787 50617 24210
rect 58031 23620 58101 24193
<< metal2 >>
rect 5532 24523 5602 24645
rect 13342 24583 13412 24655
rect 5415 24453 5602 24523
rect 13197 24513 13412 24583
rect 46613 24523 46683 24803
rect 54433 24523 54503 24738
rect 5415 24088 5485 24453
rect 13197 24091 13267 24513
rect 46528 24453 46683 24523
rect 54388 24453 54503 24523
rect 1338 19320 1408 22814
rect 9151 22643 9221 23101
rect 9151 22573 9418 22643
rect 9353 22340 9418 22573
rect 17248 22359 17318 23028
rect 17119 22289 17318 22359
rect 42407 20467 42476 24332
rect 46528 24096 46598 24453
rect 50221 22656 50291 24330
rect 54388 24089 54458 24453
rect 50221 22586 50479 22656
rect 50414 22322 50479 22586
rect 58313 22375 58383 22814
rect 58231 22305 58383 22375
<< metal3 >>
rect 19469 11839 33593 12155
rect 29059 11753 33593 11839
rect 29059 11309 32277 11753
rect 29032 9885 29260 10498
use M2_M14310591302025_256x8m81  M2_M14310591302025_256x8m81_0
timestamp 1763766357
transform 0 1 13153 -1 0 24111
box -34 -85 34 135
use M2_M14310591302025_256x8m81  M2_M14310591302025_256x8m81_1
timestamp 1763766357
transform 0 1 46496 -1 0 24100
box -34 -85 34 135
use M2_M14310591302025_256x8m81  M2_M14310591302025_256x8m81_2
timestamp 1763766357
transform 0 1 54317 -1 0 24124
box -34 -85 34 135
use M2_M14310591302025_256x8m81  M2_M14310591302025_256x8m81_3
timestamp 1763766357
transform 0 1 5426 -1 0 24122
box -34 -85 34 135
use M2_M14310591302076_256x8m81  M2_M14310591302076_256x8m81_0
timestamp 1763766357
transform -1 0 50558 0 1 23926
box -34 -281 34 281
use M2_M14310591302076_256x8m81  M2_M14310591302076_256x8m81_1
timestamp 1763766357
transform -1 0 58066 0 1 23906
box -34 -281 34 281
use M2_M14310591302076_256x8m81  M2_M14310591302076_256x8m81_2
timestamp 1763766357
transform -1 0 42748 0 1 23916
box -34 -281 34 281
use M2_M14310591302076_256x8m81  M2_M14310591302076_256x8m81_3
timestamp 1763766357
transform 1 0 9458 0 1 23928
box -34 -281 34 281
use M2_M14310591302076_256x8m81  M2_M14310591302076_256x8m81_4
timestamp 1763766357
transform 1 0 1655 0 1 23926
box -34 -281 34 281
use M2_M14310591302076_256x8m81  M2_M14310591302076_256x8m81_5
timestamp 1763766357
transform 1 0 17002 0 1 23916
box -34 -281 34 281
use M3_M24310591302077_256x8m81  M3_M24310591302077_256x8m81_0
timestamp 1763766357
transform 1 0 9141 0 1 19597
box -35 -304 35 304
use M3_M24310591302077_256x8m81  M3_M24310591302077_256x8m81_1
timestamp 1763766357
transform 1 0 17153 0 1 19603
box -35 -304 35 304
use M3_M24310591302077_256x8m81  M3_M24310591302077_256x8m81_2
timestamp 1763766357
transform 1 0 16905 0 1 19603
box -35 -304 35 304
use M3_M24310591302077_256x8m81  M3_M24310591302077_256x8m81_3
timestamp 1763766357
transform 1 0 50447 0 1 19594
box -35 -304 35 304
use M3_M24310591302077_256x8m81  M3_M24310591302077_256x8m81_4
timestamp 1763766357
transform 1 0 50202 0 1 19594
box -35 -304 35 304
use M3_M24310591302077_256x8m81  M3_M24310591302077_256x8m81_5
timestamp 1763766357
transform 1 0 58262 0 1 19593
box -35 -304 35 304
use M3_M24310591302077_256x8m81  M3_M24310591302077_256x8m81_6
timestamp 1763766357
transform 1 0 58015 0 1 19589
box -35 -304 35 304
use M3_M24310591302077_256x8m81  M3_M24310591302077_256x8m81_7
timestamp 1763766357
transform 1 0 9386 0 1 19597
box -35 -304 35 304
use M3_M24310591302078_256x8m81  M3_M24310591302078_256x8m81_0
timestamp 1763766357
transform 1 0 9141 0 1 20428
box -35 -225 35 225
use M3_M24310591302078_256x8m81  M3_M24310591302078_256x8m81_1
timestamp 1763766357
transform 1 0 17153 0 1 20434
box -35 -225 35 225
use M3_M24310591302078_256x8m81  M3_M24310591302078_256x8m81_2
timestamp 1763766357
transform 1 0 16905 0 1 20434
box -35 -225 35 225
use M3_M24310591302078_256x8m81  M3_M24310591302078_256x8m81_3
timestamp 1763766357
transform 1 0 50447 0 1 20425
box -35 -225 35 225
use M3_M24310591302078_256x8m81  M3_M24310591302078_256x8m81_4
timestamp 1763766357
transform 1 0 50202 0 1 20425
box -35 -225 35 225
use M3_M24310591302078_256x8m81  M3_M24310591302078_256x8m81_5
timestamp 1763766357
transform 1 0 58262 0 1 20424
box -35 -225 35 225
use M3_M24310591302078_256x8m81  M3_M24310591302078_256x8m81_6
timestamp 1763766357
transform 1 0 58015 0 1 20420
box -35 -225 35 225
use M3_M24310591302078_256x8m81  M3_M24310591302078_256x8m81_7
timestamp 1763766357
transform 1 0 9386 0 1 20428
box -35 -225 35 225
use M3_M24310591302079_256x8m81  M3_M24310591302079_256x8m81_0
timestamp 1763766357
transform 1 0 42441 0 1 19962
box -35 -635 35 635
use M3_M24310591302079_256x8m81  M3_M24310591302079_256x8m81_1
timestamp 1763766357
transform 1 0 1373 0 1 19972
box -35 -635 35 635
<< properties >>
string path 205.755 34.960 256.160 34.960 
<< end >>
