magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -193 28 193 46
rect -193 -28 -176 28
rect 176 -28 193 28
rect -193 -46 193 -28
<< via2 >>
rect -176 -28 176 28
<< metal3 >>
rect -193 28 193 46
rect -193 -28 -176 28
rect 176 -28 193 28
rect -193 -46 193 -28
<< end >>
