magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< polysilicon >>
rect -14 614 41 647
rect -14 -34 41 0
use nmos_5p04310591302071_512x8m81  nmos_5p04310591302071_512x8m81_0
timestamp 1763564386
transform 1 0 -14 0 1 0
box -88 -44 144 658
<< end >>
