magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< polysilicon >>
rect -42 159 13 193
rect 118 159 174 193
use pmos_5p04310591302062_3v512x8m81  pmos_5p04310591302062_3v512x8m81_0
timestamp 1763765945
transform 1 0 -14 0 1 0
box -202 -86 362 245
<< end >>
