magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
use nmos_5p04310591302084_3v1024x8m81  nmos_5p04310591302084_3v1024x8m81_0
timestamp 1764525316
transform 1 0 -14 0 1 0
box -620 -44 2662 731
<< end >>
