magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -44 181 44 198
rect -44 -161 -28 181
rect 28 -161 44 181
rect -44 -178 44 -161
<< via2 >>
rect -28 -161 28 181
<< metal3 >>
rect -45 181 45 198
rect -45 -161 -28 181
rect 28 -161 45 181
rect -45 -178 45 -161
<< end >>
