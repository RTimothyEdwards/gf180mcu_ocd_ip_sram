magic
tech gf180mcuD
magscale 1 5
timestamp 1763476864
<< metal1 >>
rect -23 124 23 133
rect -23 -124 -13 124
rect 13 -124 23 124
rect -23 -133 23 -124
<< via1 >>
rect -13 -124 13 124
<< metal2 >>
rect -23 124 23 133
rect -23 -124 -13 124
rect 13 -124 23 124
rect -23 -133 23 -124
<< end >>
