magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< polysilicon >>
rect -96 80 67 124
rect -96 52 -23 80
rect -67 -52 -23 52
rect -96 -80 -23 -52
rect 23 -80 67 80
rect -96 -124 67 -80
<< polycontact >>
rect -23 -80 23 80
<< metal1 >>
rect -39 80 39 98
rect -39 -80 -23 80
rect 23 -80 39 80
rect -39 -99 39 -80
<< end >>
