magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< metal2 >>
rect -9 190 75 215
rect -9 25 5 190
rect 61 25 75 190
rect -9 0 75 25
<< via2 >>
rect 5 25 61 190
<< metal3 >>
rect -9 190 75 215
rect -9 25 5 190
rect 61 25 75 190
rect -9 0 75 25
<< end >>
