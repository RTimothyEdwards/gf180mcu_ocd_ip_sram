VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_ocd_ip_sram__sram512x8m8wm1
  CLASS BLOCK ;
  FOREIGN gf180mcu_ocd_ip_sram__sram512x8m8wm1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 301.300 BY 329.865 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT 103.900 323.865 194.020 324.590 ;
        RECT 7.680 5.765 25.360 6.000 ;
        RECT 29.080 5.765 64.190 6.000 ;
        RECT 67.910 5.765 85.590 6.000 ;
        RECT 212.985 5.765 230.665 6.000 ;
        RECT 234.385 5.770 269.745 6.000 ;
        RECT 273.465 5.770 291.145 6.000 ;
        RECT 234.385 5.765 252.065 5.770 ;
      LAYER Metal1 ;
        RECT 4.845 319.155 5.975 319.870 ;
        RECT 4.845 318.455 6.000 319.155 ;
        RECT 295.440 318.950 296.570 319.955 ;
        RECT 295.300 318.570 296.570 318.950 ;
        RECT 4.845 317.440 5.975 318.455 ;
        RECT 295.440 317.525 296.570 318.570 ;
        RECT 4.845 313.095 5.975 313.810 ;
        RECT 4.845 312.395 6.000 313.095 ;
        RECT 295.440 312.890 296.570 313.895 ;
        RECT 295.300 312.510 296.570 312.890 ;
        RECT 4.845 311.380 5.975 312.395 ;
        RECT 295.440 311.465 296.570 312.510 ;
        RECT 4.845 307.035 5.975 307.750 ;
        RECT 4.845 306.335 6.000 307.035 ;
        RECT 295.440 306.830 296.570 307.835 ;
        RECT 295.300 306.450 296.570 306.830 ;
        RECT 4.845 305.320 5.975 306.335 ;
        RECT 295.440 305.405 296.570 306.450 ;
        RECT 4.845 300.975 5.975 301.690 ;
        RECT 4.845 300.275 6.000 300.975 ;
        RECT 295.440 300.770 296.570 301.775 ;
        RECT 295.300 300.390 296.570 300.770 ;
        RECT 4.845 299.260 5.975 300.275 ;
        RECT 295.440 299.345 296.570 300.390 ;
        RECT 4.845 294.915 5.975 295.630 ;
        RECT 4.845 294.215 6.000 294.915 ;
        RECT 295.440 294.710 296.570 295.715 ;
        RECT 295.300 294.330 296.570 294.710 ;
        RECT 4.845 293.200 5.975 294.215 ;
        RECT 295.440 293.285 296.570 294.330 ;
        RECT 4.845 288.855 5.975 289.570 ;
        RECT 4.845 288.155 6.000 288.855 ;
        RECT 295.440 288.650 296.570 289.655 ;
        RECT 295.300 288.270 296.570 288.650 ;
        RECT 4.845 287.140 5.975 288.155 ;
        RECT 295.440 287.225 296.570 288.270 ;
        RECT 4.845 282.795 5.975 283.510 ;
        RECT 4.845 282.095 6.000 282.795 ;
        RECT 295.440 282.590 296.570 283.595 ;
        RECT 295.300 282.210 296.570 282.590 ;
        RECT 4.845 281.080 5.975 282.095 ;
        RECT 295.440 281.165 296.570 282.210 ;
        RECT 4.845 276.735 5.975 277.450 ;
        RECT 4.845 276.035 6.000 276.735 ;
        RECT 295.440 276.530 296.570 277.535 ;
        RECT 295.300 276.150 296.570 276.530 ;
        RECT 4.845 275.020 5.975 276.035 ;
        RECT 295.440 275.105 296.570 276.150 ;
        RECT 4.845 270.675 5.975 271.390 ;
        RECT 4.845 269.975 6.000 270.675 ;
        RECT 295.440 270.470 296.570 271.475 ;
        RECT 295.300 270.090 296.570 270.470 ;
        RECT 4.845 268.960 5.975 269.975 ;
        RECT 295.440 269.045 296.570 270.090 ;
        RECT 4.845 264.615 5.975 265.330 ;
        RECT 4.845 263.915 6.000 264.615 ;
        RECT 295.440 264.410 296.570 265.415 ;
        RECT 295.300 264.030 296.570 264.410 ;
        RECT 4.845 262.900 5.975 263.915 ;
        RECT 295.440 262.985 296.570 264.030 ;
        RECT 4.845 258.555 5.975 259.270 ;
        RECT 4.845 257.855 6.000 258.555 ;
        RECT 295.440 258.350 296.570 259.355 ;
        RECT 295.300 257.970 296.570 258.350 ;
        RECT 4.845 256.840 5.975 257.855 ;
        RECT 295.440 256.925 296.570 257.970 ;
        RECT 4.845 252.495 5.975 253.210 ;
        RECT 4.845 251.795 6.000 252.495 ;
        RECT 295.440 252.290 296.570 253.295 ;
        RECT 295.300 251.910 296.570 252.290 ;
        RECT 4.845 250.780 5.975 251.795 ;
        RECT 295.440 250.865 296.570 251.910 ;
        RECT 4.845 246.435 5.975 247.150 ;
        RECT 4.845 245.735 6.000 246.435 ;
        RECT 295.440 246.230 296.570 247.235 ;
        RECT 295.300 245.850 296.570 246.230 ;
        RECT 4.845 244.720 5.975 245.735 ;
        RECT 295.440 244.805 296.570 245.850 ;
        RECT 4.845 240.375 5.975 241.090 ;
        RECT 4.845 239.675 6.000 240.375 ;
        RECT 295.440 240.170 296.570 241.175 ;
        RECT 295.300 239.790 296.570 240.170 ;
        RECT 4.845 238.660 5.975 239.675 ;
        RECT 295.440 238.745 296.570 239.790 ;
        RECT 4.845 234.315 5.975 235.030 ;
        RECT 4.845 233.615 6.000 234.315 ;
        RECT 295.440 234.110 296.570 235.115 ;
        RECT 295.300 233.730 296.570 234.110 ;
        RECT 4.845 232.600 5.975 233.615 ;
        RECT 295.440 232.685 296.570 233.730 ;
        RECT 4.845 228.255 5.975 228.970 ;
        RECT 4.845 227.555 6.000 228.255 ;
        RECT 295.440 228.050 296.570 229.055 ;
        RECT 295.300 227.670 296.570 228.050 ;
        RECT 4.845 226.540 5.975 227.555 ;
        RECT 295.440 226.625 296.570 227.670 ;
        RECT 4.845 222.195 5.975 222.910 ;
        RECT 4.845 221.495 6.000 222.195 ;
        RECT 295.440 221.990 296.570 222.995 ;
        RECT 295.300 221.610 296.570 221.990 ;
        RECT 4.845 220.480 5.975 221.495 ;
        RECT 295.440 220.565 296.570 221.610 ;
        RECT 4.845 216.135 5.975 216.850 ;
        RECT 4.845 215.435 6.000 216.135 ;
        RECT 295.440 215.930 296.570 216.935 ;
        RECT 295.300 215.550 296.570 215.930 ;
        RECT 4.845 214.420 5.975 215.435 ;
        RECT 295.440 214.505 296.570 215.550 ;
        RECT 4.845 210.075 5.975 210.790 ;
        RECT 4.845 209.375 6.000 210.075 ;
        RECT 295.440 209.870 296.570 210.875 ;
        RECT 295.300 209.490 296.570 209.870 ;
        RECT 4.845 208.360 5.975 209.375 ;
        RECT 295.440 208.445 296.570 209.490 ;
        RECT 4.845 204.015 5.975 204.730 ;
        RECT 4.845 203.315 6.000 204.015 ;
        RECT 295.440 203.810 296.570 204.815 ;
        RECT 295.300 203.430 296.570 203.810 ;
        RECT 4.845 202.300 5.975 203.315 ;
        RECT 295.440 202.385 296.570 203.430 ;
        RECT 4.845 197.955 5.975 198.670 ;
        RECT 4.845 197.255 6.000 197.955 ;
        RECT 295.440 197.750 296.570 198.755 ;
        RECT 295.300 197.370 296.570 197.750 ;
        RECT 4.845 196.240 5.975 197.255 ;
        RECT 295.440 196.325 296.570 197.370 ;
        RECT 4.845 191.895 5.975 192.610 ;
        RECT 4.845 191.195 6.000 191.895 ;
        RECT 295.440 191.690 296.570 192.695 ;
        RECT 295.300 191.310 296.570 191.690 ;
        RECT 4.845 190.180 5.975 191.195 ;
        RECT 295.440 190.265 296.570 191.310 ;
        RECT 4.845 185.835 5.975 186.550 ;
        RECT 4.845 185.135 6.000 185.835 ;
        RECT 295.440 185.630 296.570 186.635 ;
        RECT 295.300 185.250 296.570 185.630 ;
        RECT 4.845 184.120 5.975 185.135 ;
        RECT 295.440 184.205 296.570 185.250 ;
        RECT 4.845 179.775 5.975 180.490 ;
        RECT 4.845 179.075 6.000 179.775 ;
        RECT 295.440 179.570 296.570 180.575 ;
        RECT 295.300 179.190 296.570 179.570 ;
        RECT 4.845 178.060 5.975 179.075 ;
        RECT 295.440 178.145 296.570 179.190 ;
        RECT 4.845 173.715 5.975 174.430 ;
        RECT 4.845 173.015 6.000 173.715 ;
        RECT 295.440 173.510 296.570 174.515 ;
        RECT 295.300 173.130 296.570 173.510 ;
        RECT 4.845 172.000 5.975 173.015 ;
        RECT 295.440 172.085 296.570 173.130 ;
        RECT 4.845 167.655 5.975 168.370 ;
        RECT 4.845 166.955 6.000 167.655 ;
        RECT 295.440 167.450 296.570 168.455 ;
        RECT 295.300 167.070 296.570 167.450 ;
        RECT 4.845 165.940 5.975 166.955 ;
        RECT 295.440 166.025 296.570 167.070 ;
        RECT 4.845 161.595 5.975 162.310 ;
        RECT 4.845 160.895 6.000 161.595 ;
        RECT 295.440 161.390 296.570 162.395 ;
        RECT 295.300 161.010 296.570 161.390 ;
        RECT 4.845 159.880 5.975 160.895 ;
        RECT 295.440 159.965 296.570 161.010 ;
        RECT 4.845 155.535 5.975 156.250 ;
        RECT 4.845 154.835 6.000 155.535 ;
        RECT 295.440 155.330 296.570 156.335 ;
        RECT 295.300 154.950 296.570 155.330 ;
        RECT 4.845 153.820 5.975 154.835 ;
        RECT 295.440 153.905 296.570 154.950 ;
        RECT 4.845 149.475 5.975 150.190 ;
        RECT 4.845 148.775 6.000 149.475 ;
        RECT 295.440 149.270 296.570 150.275 ;
        RECT 295.300 148.890 296.570 149.270 ;
        RECT 4.845 147.760 5.975 148.775 ;
        RECT 295.440 147.845 296.570 148.890 ;
        RECT 4.845 143.415 5.975 144.130 ;
        RECT 4.845 142.715 6.000 143.415 ;
        RECT 295.440 143.210 296.570 144.215 ;
        RECT 295.300 142.830 296.570 143.210 ;
        RECT 4.845 141.700 5.975 142.715 ;
        RECT 295.440 141.785 296.570 142.830 ;
        RECT 4.845 137.355 5.975 138.070 ;
        RECT 4.845 136.655 6.000 137.355 ;
        RECT 295.440 137.150 296.570 138.155 ;
        RECT 295.300 136.770 296.570 137.150 ;
        RECT 4.845 135.640 5.975 136.655 ;
        RECT 295.440 135.725 296.570 136.770 ;
        RECT 4.845 131.295 5.975 132.010 ;
        RECT 4.845 130.595 6.000 131.295 ;
        RECT 295.440 131.090 296.570 132.095 ;
        RECT 295.300 130.710 296.570 131.090 ;
        RECT 4.845 129.580 5.975 130.595 ;
        RECT 295.440 129.665 296.570 130.710 ;
        RECT 4.845 125.235 5.975 125.950 ;
        RECT 4.845 124.535 6.000 125.235 ;
        RECT 295.440 125.030 296.570 126.035 ;
        RECT 295.300 124.650 296.570 125.030 ;
        RECT 4.845 123.520 5.975 124.535 ;
        RECT 295.440 123.605 296.570 124.650 ;
        RECT 93.700 5.110 95.245 6.000 ;
      LAYER Metal2 ;
        RECT 2.470 326.760 298.830 326.910 ;
        RECT 2.465 323.865 298.830 326.760 ;
        RECT 2.465 323.410 6.000 323.865 ;
        RECT 295.300 323.410 298.830 323.865 ;
        RECT 2.465 319.870 5.970 323.410 ;
        RECT 295.445 320.090 298.830 323.410 ;
        RECT 2.465 317.440 5.975 319.870 ;
        RECT 2.465 313.810 5.970 317.440 ;
        RECT 2.465 311.380 5.975 313.810 ;
        RECT 2.465 307.750 5.970 311.380 ;
        RECT 2.465 305.320 5.975 307.750 ;
        RECT 2.465 301.690 5.970 305.320 ;
        RECT 2.465 299.260 5.975 301.690 ;
        RECT 2.465 295.630 5.970 299.260 ;
        RECT 2.465 293.200 5.975 295.630 ;
        RECT 2.465 289.570 5.970 293.200 ;
        RECT 2.465 287.140 5.975 289.570 ;
        RECT 2.465 283.510 5.970 287.140 ;
        RECT 2.465 281.080 5.975 283.510 ;
        RECT 2.465 277.450 5.970 281.080 ;
        RECT 2.465 275.020 5.975 277.450 ;
        RECT 2.465 271.390 5.970 275.020 ;
        RECT 2.465 268.960 5.975 271.390 ;
        RECT 2.465 265.330 5.970 268.960 ;
        RECT 2.465 262.900 5.975 265.330 ;
        RECT 2.465 259.270 5.970 262.900 ;
        RECT 2.465 256.840 5.975 259.270 ;
        RECT 2.465 253.210 5.970 256.840 ;
        RECT 2.465 250.780 5.975 253.210 ;
        RECT 2.465 247.150 5.970 250.780 ;
        RECT 2.465 244.720 5.975 247.150 ;
        RECT 2.465 241.090 5.970 244.720 ;
        RECT 2.465 238.660 5.975 241.090 ;
        RECT 2.465 235.030 5.970 238.660 ;
        RECT 2.465 232.600 5.975 235.030 ;
        RECT 2.465 228.970 5.970 232.600 ;
        RECT 2.465 226.540 5.975 228.970 ;
        RECT 2.465 222.910 5.970 226.540 ;
        RECT 2.465 220.480 5.975 222.910 ;
        RECT 2.465 216.850 5.970 220.480 ;
        RECT 2.465 214.420 5.975 216.850 ;
        RECT 2.465 210.790 5.970 214.420 ;
        RECT 2.465 208.360 5.975 210.790 ;
        RECT 2.465 204.730 5.970 208.360 ;
        RECT 2.465 202.300 5.975 204.730 ;
        RECT 2.465 198.670 5.970 202.300 ;
        RECT 2.465 196.240 5.975 198.670 ;
        RECT 2.465 192.610 5.970 196.240 ;
        RECT 2.465 190.180 5.975 192.610 ;
        RECT 2.465 186.550 5.970 190.180 ;
        RECT 2.465 184.120 5.975 186.550 ;
        RECT 2.465 180.490 5.970 184.120 ;
        RECT 2.465 178.060 5.975 180.490 ;
        RECT 2.465 174.430 5.970 178.060 ;
        RECT 295.440 176.180 298.830 320.090 ;
        RECT 2.465 172.000 5.975 174.430 ;
        RECT 2.465 168.370 5.970 172.000 ;
        RECT 2.465 165.940 5.975 168.370 ;
        RECT 2.465 162.310 5.970 165.940 ;
        RECT 2.465 159.880 5.975 162.310 ;
        RECT 2.465 156.250 5.970 159.880 ;
        RECT 2.465 153.820 5.975 156.250 ;
        RECT 2.465 150.190 5.970 153.820 ;
        RECT 2.465 147.760 5.975 150.190 ;
        RECT 2.465 144.130 5.970 147.760 ;
        RECT 2.465 141.700 5.975 144.130 ;
        RECT 2.465 138.070 5.970 141.700 ;
        RECT 2.465 135.640 5.975 138.070 ;
        RECT 2.465 132.010 5.970 135.640 ;
        RECT 2.465 129.580 5.975 132.010 ;
        RECT 2.465 125.950 5.970 129.580 ;
        RECT 2.465 123.520 5.975 125.950 ;
        RECT 2.465 118.255 5.970 123.520 ;
        RECT 295.440 118.255 298.835 176.180 ;
        RECT 2.465 41.740 5.975 118.255 ;
        RECT 295.330 41.740 298.835 118.255 ;
        RECT 2.465 39.990 5.970 41.740 ;
        RECT 295.330 39.990 298.830 41.740 ;
        RECT 2.465 1.410 5.975 39.990 ;
        RECT 26.795 4.830 27.580 6.000 ;
        RECT 65.605 4.830 66.390 6.000 ;
        RECT 88.750 4.310 89.535 6.000 ;
        RECT 93.695 5.965 95.245 6.000 ;
        RECT 131.250 5.180 132.035 6.000 ;
        RECT 137.620 5.180 138.405 6.000 ;
        RECT 202.670 4.505 204.220 6.000 ;
        RECT 207.850 4.310 208.635 6.000 ;
        RECT 232.070 4.830 232.855 6.000 ;
        RECT 271.220 4.830 272.005 6.000 ;
        RECT 2.470 0.985 5.975 1.410 ;
        RECT 295.330 0.985 298.835 39.990 ;
        RECT 2.475 0.980 5.975 0.985 ;
        RECT 295.335 0.980 298.835 0.985 ;
      LAYER Metal3 ;
        RECT 5.050 329.705 8.550 329.710 ;
        RECT 5.050 327.580 8.555 329.705 ;
        RECT 14.475 327.580 17.975 329.710 ;
        RECT 24.600 329.705 28.100 329.710 ;
        RECT 24.600 327.580 28.105 329.705 ;
        RECT 33.375 327.580 36.875 329.710 ;
        RECT 44.150 329.705 47.650 329.710 ;
        RECT 44.150 327.580 47.655 329.705 ;
        RECT 52.275 327.580 55.775 329.710 ;
        RECT 63.700 329.705 67.200 329.710 ;
        RECT 63.700 327.580 67.205 329.705 ;
        RECT 5.060 326.910 8.555 327.580 ;
        RECT 14.480 326.910 17.975 327.580 ;
        RECT 24.610 326.910 28.105 327.580 ;
        RECT 33.380 326.910 36.875 327.580 ;
        RECT 44.160 326.910 47.655 327.580 ;
        RECT 52.280 326.910 55.775 327.580 ;
        RECT 63.710 326.910 67.205 327.580 ;
        RECT 72.285 327.580 75.785 329.710 ;
        RECT 84.740 327.580 88.240 329.710 ;
        RECT 72.285 326.910 75.780 327.580 ;
        RECT 84.745 326.910 88.240 327.580 ;
        RECT 93.000 327.580 96.500 329.710 ;
        RECT 107.485 327.580 110.985 329.710 ;
        RECT 123.950 327.580 127.450 329.710 ;
        RECT 135.045 327.580 138.545 329.710 ;
        RECT 144.305 327.580 147.805 329.710 ;
        RECT 157.740 327.580 161.240 329.710 ;
        RECT 162.095 327.580 165.595 329.710 ;
        RECT 171.150 327.580 174.650 329.710 ;
        RECT 93.000 326.910 96.495 327.580 ;
        RECT 107.485 326.910 110.980 327.580 ;
        RECT 123.950 326.910 127.445 327.580 ;
        RECT 135.045 326.910 138.540 327.580 ;
        RECT 144.305 326.910 147.800 327.580 ;
        RECT 157.740 326.910 161.235 327.580 ;
        RECT 162.095 326.910 165.590 327.580 ;
        RECT 171.155 326.910 174.650 327.580 ;
        RECT 183.990 327.580 187.490 329.710 ;
        RECT 189.915 327.580 193.415 329.710 ;
        RECT 201.410 328.095 204.910 329.710 ;
        RECT 210.515 329.705 214.015 329.710 ;
        RECT 210.515 328.240 214.020 329.705 ;
        RECT 183.990 326.910 187.485 327.580 ;
        RECT 189.915 326.910 193.410 327.580 ;
        RECT 201.415 326.910 204.910 328.095 ;
        RECT 210.510 327.575 214.020 328.240 ;
        RECT 210.525 326.910 214.020 327.575 ;
        RECT 221.995 327.580 225.495 329.710 ;
        RECT 230.065 327.580 233.565 329.710 ;
        RECT 240.895 327.580 244.395 329.710 ;
        RECT 249.565 329.705 253.065 329.710 ;
        RECT 249.565 327.580 253.070 329.705 ;
        RECT 221.995 326.910 225.490 327.580 ;
        RECT 230.065 326.910 233.560 327.580 ;
        RECT 240.895 326.910 244.390 327.580 ;
        RECT 249.575 326.910 253.070 327.580 ;
        RECT 259.795 327.580 263.295 329.710 ;
        RECT 269.115 329.705 272.615 329.710 ;
        RECT 269.115 327.580 272.620 329.705 ;
        RECT 259.795 326.910 263.290 327.580 ;
        RECT 269.125 326.910 272.620 327.580 ;
        RECT 279.300 327.580 282.800 329.710 ;
        RECT 290.105 327.580 293.605 329.710 ;
        RECT 279.300 326.910 282.795 327.580 ;
        RECT 290.110 326.910 293.605 327.580 ;
        RECT 295.330 327.580 298.830 329.710 ;
        RECT 295.330 326.910 298.825 327.580 ;
        RECT 0.000 323.865 301.300 326.910 ;
        RECT 0.000 323.410 6.000 323.865 ;
        RECT 295.300 323.410 301.300 323.865 ;
        RECT 5.060 323.405 6.000 323.410 ;
        RECT 296.440 319.955 301.300 319.965 ;
        RECT 0.000 317.430 5.975 319.880 ;
        RECT 295.440 317.525 301.300 319.955 ;
        RECT 296.440 317.515 301.300 317.525 ;
        RECT 296.440 313.895 301.300 313.905 ;
        RECT 0.000 311.370 5.975 313.820 ;
        RECT 295.440 311.465 301.300 313.895 ;
        RECT 296.440 311.455 301.300 311.465 ;
        RECT 296.440 307.835 301.300 307.845 ;
        RECT 0.000 305.310 5.975 307.760 ;
        RECT 295.440 305.405 301.300 307.835 ;
        RECT 296.440 305.395 301.300 305.405 ;
        RECT 296.440 301.775 301.300 301.785 ;
        RECT 0.000 299.250 5.975 301.700 ;
        RECT 295.440 299.345 301.300 301.775 ;
        RECT 296.440 299.335 301.300 299.345 ;
        RECT 296.440 295.715 301.300 295.725 ;
        RECT 0.000 293.190 5.975 295.640 ;
        RECT 295.440 293.285 301.300 295.715 ;
        RECT 296.440 293.275 301.300 293.285 ;
        RECT 296.440 289.655 301.300 289.665 ;
        RECT 0.000 287.130 5.975 289.580 ;
        RECT 295.440 287.225 301.300 289.655 ;
        RECT 296.440 287.215 301.300 287.225 ;
        RECT 296.440 283.595 301.300 283.605 ;
        RECT 0.000 281.070 5.975 283.520 ;
        RECT 295.440 281.165 301.300 283.595 ;
        RECT 296.440 281.155 301.300 281.165 ;
        RECT 296.440 277.535 301.300 277.545 ;
        RECT 0.000 275.010 5.975 277.460 ;
        RECT 295.440 275.105 301.300 277.535 ;
        RECT 296.440 275.095 301.300 275.105 ;
        RECT 296.440 271.475 301.300 271.485 ;
        RECT 0.000 268.950 5.975 271.400 ;
        RECT 295.440 269.045 301.300 271.475 ;
        RECT 296.440 269.035 301.300 269.045 ;
        RECT 296.440 265.415 301.300 265.425 ;
        RECT 0.000 262.890 5.975 265.340 ;
        RECT 295.440 262.985 301.300 265.415 ;
        RECT 296.440 262.975 301.300 262.985 ;
        RECT 296.440 259.355 301.300 259.365 ;
        RECT 0.000 256.830 5.975 259.280 ;
        RECT 295.440 256.925 301.300 259.355 ;
        RECT 296.440 256.915 301.300 256.925 ;
        RECT 296.440 253.295 301.300 253.305 ;
        RECT 0.000 250.770 5.975 253.220 ;
        RECT 295.440 250.865 301.300 253.295 ;
        RECT 296.440 250.855 301.300 250.865 ;
        RECT 296.440 247.235 301.300 247.245 ;
        RECT 0.000 244.710 5.975 247.160 ;
        RECT 295.440 244.805 301.300 247.235 ;
        RECT 296.440 244.795 301.300 244.805 ;
        RECT 296.440 241.175 301.300 241.185 ;
        RECT 0.000 238.650 5.975 241.100 ;
        RECT 295.440 238.745 301.300 241.175 ;
        RECT 296.440 238.735 301.300 238.745 ;
        RECT 296.440 235.115 301.300 235.125 ;
        RECT 0.000 232.590 5.975 235.040 ;
        RECT 295.440 232.685 301.300 235.115 ;
        RECT 296.440 232.675 301.300 232.685 ;
        RECT 296.440 229.055 301.300 229.065 ;
        RECT 0.000 226.530 5.975 228.980 ;
        RECT 295.440 226.625 301.300 229.055 ;
        RECT 296.440 226.615 301.300 226.625 ;
        RECT 296.440 222.995 301.300 223.005 ;
        RECT 0.000 220.470 5.975 222.920 ;
        RECT 295.440 220.565 301.300 222.995 ;
        RECT 296.440 220.555 301.300 220.565 ;
        RECT 296.440 216.935 301.300 216.945 ;
        RECT 0.000 214.410 5.975 216.860 ;
        RECT 295.440 214.505 301.300 216.935 ;
        RECT 296.440 214.495 301.300 214.505 ;
        RECT 296.440 210.875 301.300 210.885 ;
        RECT 0.000 208.350 5.975 210.800 ;
        RECT 295.440 208.445 301.300 210.875 ;
        RECT 296.440 208.435 301.300 208.445 ;
        RECT 296.440 204.815 301.300 204.825 ;
        RECT 0.000 202.290 5.975 204.740 ;
        RECT 295.440 202.385 301.300 204.815 ;
        RECT 296.440 202.375 301.300 202.385 ;
        RECT 296.440 198.755 301.300 198.765 ;
        RECT 0.000 196.230 5.975 198.680 ;
        RECT 295.440 196.325 301.300 198.755 ;
        RECT 296.440 196.315 301.300 196.325 ;
        RECT 296.440 192.695 301.300 192.705 ;
        RECT 0.000 190.170 5.975 192.620 ;
        RECT 295.440 190.265 301.300 192.695 ;
        RECT 296.440 190.255 301.300 190.265 ;
        RECT 296.440 186.635 301.300 186.645 ;
        RECT 0.000 184.110 5.975 186.560 ;
        RECT 295.440 184.205 301.300 186.635 ;
        RECT 296.440 184.195 301.300 184.205 ;
        RECT 296.440 180.575 301.300 180.585 ;
        RECT 0.000 178.050 5.975 180.500 ;
        RECT 295.440 178.145 301.300 180.575 ;
        RECT 296.440 178.135 301.300 178.145 ;
        RECT 296.440 174.515 301.300 174.525 ;
        RECT 0.000 171.990 5.975 174.440 ;
        RECT 295.440 172.085 301.300 174.515 ;
        RECT 296.440 172.075 301.300 172.085 ;
        RECT 296.440 168.455 301.300 168.465 ;
        RECT 0.000 165.930 5.975 168.380 ;
        RECT 295.440 166.025 301.300 168.455 ;
        RECT 296.440 166.015 301.300 166.025 ;
        RECT 296.440 162.395 301.300 162.405 ;
        RECT 0.000 159.870 5.975 162.320 ;
        RECT 295.440 159.965 301.300 162.395 ;
        RECT 296.440 159.955 301.300 159.965 ;
        RECT 296.440 156.335 301.300 156.345 ;
        RECT 0.000 153.810 5.975 156.260 ;
        RECT 295.440 153.905 301.300 156.335 ;
        RECT 296.440 153.895 301.300 153.905 ;
        RECT 296.440 150.275 301.300 150.285 ;
        RECT 0.000 147.750 5.975 150.200 ;
        RECT 295.440 147.845 301.300 150.275 ;
        RECT 296.440 147.835 301.300 147.845 ;
        RECT 296.440 144.215 301.300 144.225 ;
        RECT 0.000 141.690 5.975 144.140 ;
        RECT 295.440 141.785 301.300 144.215 ;
        RECT 296.440 141.775 301.300 141.785 ;
        RECT 296.440 138.155 301.300 138.165 ;
        RECT 0.000 135.630 5.975 138.080 ;
        RECT 295.440 135.725 301.300 138.155 ;
        RECT 296.440 135.715 301.300 135.725 ;
        RECT 296.440 132.095 301.300 132.105 ;
        RECT 0.000 129.570 5.975 132.020 ;
        RECT 295.440 129.665 301.300 132.095 ;
        RECT 296.440 129.655 301.300 129.665 ;
        RECT 296.440 126.035 301.300 126.045 ;
        RECT 0.000 123.510 5.975 125.960 ;
        RECT 295.440 123.605 301.300 126.035 ;
        RECT 296.440 123.595 301.300 123.605 ;
        RECT 0.000 117.725 3.545 117.730 ;
        RECT 297.750 117.725 301.300 117.730 ;
        RECT 0.000 110.700 6.000 117.725 ;
        RECT 295.300 110.700 301.300 117.725 ;
        RECT 0.000 103.990 5.975 110.700 ;
        RECT 295.335 103.990 301.300 110.700 ;
        RECT 0.000 102.995 6.000 103.990 ;
        RECT 295.300 102.995 301.300 103.990 ;
        RECT 300.600 102.990 301.300 102.995 ;
        RECT 0.000 84.070 3.545 84.075 ;
        RECT 297.750 84.070 301.300 84.075 ;
        RECT 0.000 82.120 5.975 84.070 ;
        RECT 295.335 82.120 301.300 84.070 ;
        RECT 0.000 80.575 6.000 82.120 ;
        RECT 0.010 80.570 6.000 80.575 ;
        RECT 295.300 80.570 301.300 82.120 ;
        RECT 0.000 72.575 3.545 72.630 ;
        RECT 297.750 72.575 301.300 72.580 ;
        RECT 0.000 63.100 6.000 72.575 ;
        RECT 0.010 63.045 6.000 63.100 ;
        RECT 295.300 63.045 301.300 72.575 ;
        RECT 0.000 49.610 3.545 49.665 ;
        RECT 297.750 49.610 301.300 49.615 ;
        RECT 0.000 47.105 6.000 49.610 ;
        RECT 295.300 47.105 301.300 49.610 ;
        RECT 0.000 44.950 5.975 47.105 ;
        RECT 295.335 44.950 301.300 47.105 ;
        RECT 0.000 42.170 6.000 44.950 ;
        RECT 0.010 42.115 6.000 42.170 ;
        RECT 295.300 42.115 301.300 44.950 ;
        RECT 0.000 33.290 3.545 33.345 ;
        RECT 297.750 33.290 301.300 33.295 ;
        RECT 0.000 28.575 6.000 33.290 ;
        RECT 0.010 28.520 6.000 28.575 ;
        RECT 295.300 28.520 301.300 33.290 ;
        RECT 0.000 19.730 3.545 19.745 ;
        RECT 0.000 19.690 5.915 19.730 ;
        RECT 295.395 19.695 298.695 19.730 ;
        RECT 0.000 18.095 6.000 19.690 ;
        RECT 295.300 18.095 301.300 19.695 ;
        RECT 0.000 15.790 5.995 18.095 ;
        RECT 295.315 15.800 301.300 18.095 ;
        RECT 0.000 14.255 6.000 15.790 ;
        RECT 0.010 14.200 6.000 14.255 ;
        RECT 295.300 14.200 301.300 15.800 ;
        RECT 0.000 6.000 6.000 7.810 ;
        RECT 295.330 7.805 301.300 7.810 ;
        RECT 295.300 6.000 301.300 7.805 ;
        RECT 0.000 4.310 301.300 6.000 ;
        RECT 0.010 4.305 10.635 4.310 ;
        RECT 2.465 0.000 5.970 4.305 ;
        RECT 7.135 0.000 10.635 4.305 ;
        RECT 12.045 0.000 15.545 4.310 ;
        RECT 20.445 0.000 23.945 4.310 ;
        RECT 24.645 0.000 28.145 4.310 ;
        RECT 28.845 0.000 32.345 4.310 ;
        RECT 37.245 0.000 40.745 4.310 ;
        RECT 43.550 0.000 47.050 4.310 ;
        RECT 49.845 0.000 53.345 4.310 ;
        RECT 58.245 0.000 61.745 4.310 ;
        RECT 62.445 0.000 65.945 4.310 ;
        RECT 66.645 0.000 70.145 4.310 ;
        RECT 76.685 0.000 80.185 4.310 ;
        RECT 80.885 0.000 84.385 4.310 ;
        RECT 85.435 0.000 88.935 4.310 ;
        RECT 89.985 0.000 93.485 4.310 ;
        RECT 94.535 0.000 98.035 4.310 ;
        RECT 99.085 0.000 102.585 4.310 ;
        RECT 103.635 0.000 107.135 4.310 ;
        RECT 126.105 0.000 129.605 4.310 ;
        RECT 137.295 0.000 140.795 4.310 ;
        RECT 148.515 0.000 152.015 4.310 ;
        RECT 156.915 0.000 160.415 4.310 ;
        RECT 165.315 0.000 168.815 4.310 ;
        RECT 169.980 0.000 173.480 4.310 ;
        RECT 174.565 0.000 178.065 4.310 ;
        RECT 190.600 0.000 194.100 4.310 ;
        RECT 195.150 0.000 198.650 4.310 ;
        RECT 199.700 0.000 203.200 4.310 ;
        RECT 204.250 0.000 207.750 4.310 ;
        RECT 208.800 0.000 212.300 4.310 ;
        RECT 213.350 0.000 216.850 4.310 ;
        RECT 218.030 0.000 221.530 4.310 ;
        RECT 227.960 0.000 231.460 4.310 ;
        RECT 232.160 0.000 235.660 4.310 ;
        RECT 236.360 0.000 239.860 4.310 ;
        RECT 244.760 0.000 248.260 4.310 ;
        RECT 251.055 0.000 254.555 4.310 ;
        RECT 257.360 0.000 260.860 4.310 ;
        RECT 265.760 0.000 269.260 4.310 ;
        RECT 269.960 0.000 273.460 4.310 ;
        RECT 274.160 0.000 277.660 4.310 ;
        RECT 283.560 0.000 287.060 4.310 ;
        RECT 288.465 4.305 301.300 4.310 ;
        RECT 288.465 0.000 291.965 4.305 ;
        RECT 295.330 0.000 298.830 4.305 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.985 325.185 300.315 328.720 ;
        RECT 0.985 322.855 4.485 325.185 ;
        RECT 7.360 323.865 7.935 325.185 ;
        RECT 26.910 323.865 27.485 325.185 ;
        RECT 46.460 323.865 47.035 325.185 ;
        RECT 66.010 323.865 66.585 325.185 ;
        RECT 85.365 323.865 85.940 325.185 ;
        RECT 90.140 323.865 92.685 325.185 ;
        RECT 96.620 324.850 102.185 325.185 ;
        RECT 95.855 323.865 102.185 324.850 ;
        RECT 119.790 323.865 122.545 325.185 ;
        RECT 140.215 323.865 142.065 325.185 ;
        RECT 153.080 323.865 155.970 325.185 ;
        RECT 175.340 323.865 178.195 325.185 ;
        RECT 194.845 323.865 202.075 325.185 ;
        RECT 204.765 323.865 207.310 325.185 ;
        RECT 212.825 323.865 213.400 325.185 ;
        RECT 232.365 323.865 232.940 325.185 ;
        RECT 251.875 323.865 252.450 325.185 ;
        RECT 271.425 323.865 272.000 325.185 ;
        RECT 290.730 323.865 291.305 325.185 ;
        RECT 296.815 323.005 300.315 325.185 ;
        RECT 0.985 322.705 4.490 322.855 ;
        RECT 0.985 320.900 6.000 322.705 ;
        RECT 0.985 317.605 4.490 320.900 ;
        RECT 296.815 320.575 301.300 323.005 ;
        RECT 0.985 316.795 4.485 317.605 ;
        RECT 296.815 316.945 300.315 320.575 ;
        RECT 0.985 316.645 4.490 316.795 ;
        RECT 0.985 314.840 6.000 316.645 ;
        RECT 0.985 311.545 4.490 314.840 ;
        RECT 296.815 314.515 301.300 316.945 ;
        RECT 0.985 310.735 4.485 311.545 ;
        RECT 296.815 310.885 300.315 314.515 ;
        RECT 0.985 310.585 4.490 310.735 ;
        RECT 0.985 308.780 6.000 310.585 ;
        RECT 0.985 305.485 4.490 308.780 ;
        RECT 296.815 308.455 301.300 310.885 ;
        RECT 0.985 304.675 4.485 305.485 ;
        RECT 296.815 304.825 300.315 308.455 ;
        RECT 0.985 304.525 4.490 304.675 ;
        RECT 0.985 302.720 6.000 304.525 ;
        RECT 0.985 299.425 4.490 302.720 ;
        RECT 296.815 302.395 301.300 304.825 ;
        RECT 0.985 298.615 4.485 299.425 ;
        RECT 296.815 298.765 300.315 302.395 ;
        RECT 0.985 298.465 4.490 298.615 ;
        RECT 0.985 296.660 6.000 298.465 ;
        RECT 295.300 297.230 296.325 297.930 ;
        RECT 0.985 293.365 4.490 296.660 ;
        RECT 296.815 296.335 301.300 298.765 ;
        RECT 0.985 292.555 4.485 293.365 ;
        RECT 296.815 292.705 300.315 296.335 ;
        RECT 0.985 292.405 4.490 292.555 ;
        RECT 0.985 290.600 6.000 292.405 ;
        RECT 0.985 287.305 4.490 290.600 ;
        RECT 296.815 290.275 301.300 292.705 ;
        RECT 0.985 286.495 4.485 287.305 ;
        RECT 296.815 286.645 300.315 290.275 ;
        RECT 0.985 286.345 4.490 286.495 ;
        RECT 0.985 284.540 6.000 286.345 ;
        RECT 0.985 281.245 4.490 284.540 ;
        RECT 296.815 284.215 301.300 286.645 ;
        RECT 0.985 280.435 4.485 281.245 ;
        RECT 296.815 280.585 300.315 284.215 ;
        RECT 0.985 280.285 4.490 280.435 ;
        RECT 0.985 278.480 6.000 280.285 ;
        RECT 0.985 275.185 4.490 278.480 ;
        RECT 296.815 278.155 301.300 280.585 ;
        RECT 0.985 274.375 4.485 275.185 ;
        RECT 296.815 274.525 300.315 278.155 ;
        RECT 0.985 274.225 4.490 274.375 ;
        RECT 0.985 272.420 6.000 274.225 ;
        RECT 0.985 269.125 4.490 272.420 ;
        RECT 296.815 272.095 301.300 274.525 ;
        RECT 0.985 268.315 4.485 269.125 ;
        RECT 296.815 268.465 300.315 272.095 ;
        RECT 0.985 268.165 4.490 268.315 ;
        RECT 0.985 266.360 6.000 268.165 ;
        RECT 0.985 263.065 4.490 266.360 ;
        RECT 296.815 266.035 301.300 268.465 ;
        RECT 0.985 262.255 4.485 263.065 ;
        RECT 296.815 262.405 300.315 266.035 ;
        RECT 0.985 262.105 4.490 262.255 ;
        RECT 0.985 260.300 6.000 262.105 ;
        RECT 0.985 257.005 4.490 260.300 ;
        RECT 296.815 259.975 301.300 262.405 ;
        RECT 0.985 256.195 4.485 257.005 ;
        RECT 296.815 256.345 300.315 259.975 ;
        RECT 0.985 256.045 4.490 256.195 ;
        RECT 0.985 254.240 6.000 256.045 ;
        RECT 0.985 250.945 4.490 254.240 ;
        RECT 296.815 253.915 301.300 256.345 ;
        RECT 0.985 250.135 4.485 250.945 ;
        RECT 296.815 250.285 300.315 253.915 ;
        RECT 0.985 249.985 4.490 250.135 ;
        RECT 0.985 248.180 6.000 249.985 ;
        RECT 0.985 244.885 4.490 248.180 ;
        RECT 296.815 247.855 301.300 250.285 ;
        RECT 0.985 244.075 4.485 244.885 ;
        RECT 296.815 244.225 300.315 247.855 ;
        RECT 0.985 243.925 4.490 244.075 ;
        RECT 0.985 242.120 6.000 243.925 ;
        RECT 0.985 238.825 4.490 242.120 ;
        RECT 296.815 241.795 301.300 244.225 ;
        RECT 0.985 238.015 4.485 238.825 ;
        RECT 296.815 238.165 300.315 241.795 ;
        RECT 0.985 237.865 4.490 238.015 ;
        RECT 0.985 236.060 6.000 237.865 ;
        RECT 0.985 232.765 4.490 236.060 ;
        RECT 296.815 235.735 301.300 238.165 ;
        RECT 0.985 231.955 4.485 232.765 ;
        RECT 296.815 232.105 300.315 235.735 ;
        RECT 0.985 231.805 4.490 231.955 ;
        RECT 0.985 230.000 6.000 231.805 ;
        RECT 0.985 226.705 4.490 230.000 ;
        RECT 296.815 229.675 301.300 232.105 ;
        RECT 0.985 225.895 4.485 226.705 ;
        RECT 296.815 226.045 300.315 229.675 ;
        RECT 0.985 225.745 4.490 225.895 ;
        RECT 0.985 223.940 6.000 225.745 ;
        RECT 0.985 220.645 4.490 223.940 ;
        RECT 296.815 223.615 301.300 226.045 ;
        RECT 0.985 219.835 4.485 220.645 ;
        RECT 296.815 219.985 300.315 223.615 ;
        RECT 0.985 219.685 4.490 219.835 ;
        RECT 0.985 217.880 6.000 219.685 ;
        RECT 0.985 214.585 4.490 217.880 ;
        RECT 296.815 217.555 301.300 219.985 ;
        RECT 0.985 213.775 4.485 214.585 ;
        RECT 296.815 213.925 300.315 217.555 ;
        RECT 0.985 213.625 4.490 213.775 ;
        RECT 0.985 211.820 6.000 213.625 ;
        RECT 0.985 208.525 4.490 211.820 ;
        RECT 296.815 211.495 301.300 213.925 ;
        RECT 0.985 207.715 4.485 208.525 ;
        RECT 296.815 207.865 300.315 211.495 ;
        RECT 0.985 207.565 4.490 207.715 ;
        RECT 0.985 205.760 6.000 207.565 ;
        RECT 0.985 202.465 4.490 205.760 ;
        RECT 296.815 205.435 301.300 207.865 ;
        RECT 0.985 201.655 4.485 202.465 ;
        RECT 296.815 201.805 300.315 205.435 ;
        RECT 0.985 201.505 4.490 201.655 ;
        RECT 0.985 199.700 6.000 201.505 ;
        RECT 0.985 196.405 4.490 199.700 ;
        RECT 296.815 199.375 301.300 201.805 ;
        RECT 0.985 195.595 4.485 196.405 ;
        RECT 296.815 195.745 300.315 199.375 ;
        RECT 0.985 195.445 4.490 195.595 ;
        RECT 0.985 193.640 6.000 195.445 ;
        RECT 0.985 190.345 4.490 193.640 ;
        RECT 296.815 193.315 301.300 195.745 ;
        RECT 0.985 189.535 4.485 190.345 ;
        RECT 296.815 189.685 300.315 193.315 ;
        RECT 0.985 189.385 4.490 189.535 ;
        RECT 0.985 187.580 6.000 189.385 ;
        RECT 0.985 184.285 4.490 187.580 ;
        RECT 296.815 187.255 301.300 189.685 ;
        RECT 0.985 183.475 4.485 184.285 ;
        RECT 296.815 183.625 300.315 187.255 ;
        RECT 0.985 183.325 4.490 183.475 ;
        RECT 0.985 181.520 6.000 183.325 ;
        RECT 0.985 178.225 4.490 181.520 ;
        RECT 296.815 181.195 301.300 183.625 ;
        RECT 0.985 177.415 4.485 178.225 ;
        RECT 296.815 177.565 300.315 181.195 ;
        RECT 0.985 177.265 4.490 177.415 ;
        RECT 0.985 175.460 6.000 177.265 ;
        RECT 0.985 172.165 4.490 175.460 ;
        RECT 296.815 175.135 301.300 177.565 ;
        RECT 0.985 171.355 4.485 172.165 ;
        RECT 296.815 171.505 300.315 175.135 ;
        RECT 0.985 171.205 4.490 171.355 ;
        RECT 0.985 169.400 6.000 171.205 ;
        RECT 0.985 166.105 4.490 169.400 ;
        RECT 296.815 169.075 301.300 171.505 ;
        RECT 0.985 165.295 4.485 166.105 ;
        RECT 296.815 165.445 300.315 169.075 ;
        RECT 0.985 165.145 4.490 165.295 ;
        RECT 0.985 163.340 6.000 165.145 ;
        RECT 0.985 160.045 4.490 163.340 ;
        RECT 296.815 163.015 301.300 165.445 ;
        RECT 0.985 159.235 4.485 160.045 ;
        RECT 296.815 159.385 300.315 163.015 ;
        RECT 0.985 159.085 4.490 159.235 ;
        RECT 0.985 157.280 6.000 159.085 ;
        RECT 0.985 153.985 4.490 157.280 ;
        RECT 296.815 156.955 301.300 159.385 ;
        RECT 0.985 153.175 4.485 153.985 ;
        RECT 296.815 153.325 300.315 156.955 ;
        RECT 0.985 153.025 4.490 153.175 ;
        RECT 0.985 151.220 6.000 153.025 ;
        RECT 0.985 147.925 4.490 151.220 ;
        RECT 296.815 150.895 301.300 153.325 ;
        RECT 0.985 147.115 4.485 147.925 ;
        RECT 296.815 147.265 300.315 150.895 ;
        RECT 0.985 146.965 4.490 147.115 ;
        RECT 0.985 145.160 6.000 146.965 ;
        RECT 0.985 141.865 4.490 145.160 ;
        RECT 296.815 144.835 301.300 147.265 ;
        RECT 0.985 141.055 4.485 141.865 ;
        RECT 296.815 141.205 300.315 144.835 ;
        RECT 0.985 140.905 4.490 141.055 ;
        RECT 0.985 139.100 6.000 140.905 ;
        RECT 0.985 135.805 4.490 139.100 ;
        RECT 296.815 138.775 301.300 141.205 ;
        RECT 0.985 134.995 4.485 135.805 ;
        RECT 296.815 135.145 300.315 138.775 ;
        RECT 0.985 134.845 4.490 134.995 ;
        RECT 0.985 133.040 6.000 134.845 ;
        RECT 0.985 129.745 4.490 133.040 ;
        RECT 296.815 132.715 301.300 135.145 ;
        RECT 0.985 128.935 4.485 129.745 ;
        RECT 296.815 129.085 300.315 132.715 ;
        RECT 0.985 128.785 4.490 128.935 ;
        RECT 0.985 126.980 6.000 128.785 ;
        RECT 0.985 123.685 4.490 126.980 ;
        RECT 296.815 126.655 301.300 129.085 ;
        RECT 0.985 95.085 4.485 123.685 ;
        RECT 296.815 122.785 300.315 126.655 ;
        RECT 295.300 122.175 300.315 122.785 ;
        RECT 296.815 120.225 300.315 122.175 ;
        RECT 295.300 119.630 300.315 120.225 ;
        RECT 296.815 95.085 300.315 119.630 ;
        RECT 0.985 94.615 6.000 95.085 ;
        RECT 295.300 94.615 300.315 95.085 ;
        RECT 0.985 77.060 4.485 94.615 ;
        RECT 296.815 77.060 300.315 94.615 ;
        RECT 0.985 76.380 6.000 77.060 ;
        RECT 295.300 76.380 300.315 77.060 ;
        RECT 0.985 4.485 4.485 76.380 ;
        RECT 95.850 5.030 97.395 6.000 ;
        RECT 100.195 5.030 140.625 6.000 ;
        RECT 177.920 5.030 198.050 6.000 ;
        RECT 200.530 5.030 202.075 6.000 ;
        RECT 95.850 4.485 202.075 5.030 ;
        RECT 296.815 4.485 300.315 76.380 ;
        RECT 0.985 0.985 300.315 4.485 ;
      LAYER Metal2 ;
        RECT 0.985 327.580 300.315 328.720 ;
        RECT 0.995 320.590 2.125 323.020 ;
        RECT 300.170 320.575 301.300 323.005 ;
        RECT 0.995 314.530 2.125 316.960 ;
        RECT 300.170 314.515 301.300 316.945 ;
        RECT 0.995 308.470 2.125 310.900 ;
        RECT 300.170 308.455 301.300 310.885 ;
        RECT 0.995 302.410 2.125 304.840 ;
        RECT 300.170 302.395 301.300 304.825 ;
        RECT 0.995 296.350 2.125 298.780 ;
        RECT 300.170 296.335 301.300 298.765 ;
        RECT 0.995 290.290 2.125 292.720 ;
        RECT 300.170 290.275 301.300 292.705 ;
        RECT 0.995 284.230 2.125 286.660 ;
        RECT 300.170 284.215 301.300 286.645 ;
        RECT 0.995 278.170 2.125 280.600 ;
        RECT 300.170 278.155 301.300 280.585 ;
        RECT 0.995 272.110 2.125 274.540 ;
        RECT 300.170 272.095 301.300 274.525 ;
        RECT 0.995 266.050 2.125 268.480 ;
        RECT 300.170 266.035 301.300 268.465 ;
        RECT 0.995 259.990 2.125 262.420 ;
        RECT 300.170 259.975 301.300 262.405 ;
        RECT 0.995 253.930 2.125 256.360 ;
        RECT 300.170 253.915 301.300 256.345 ;
        RECT 0.995 247.870 2.125 250.300 ;
        RECT 300.170 247.855 301.300 250.285 ;
        RECT 0.995 241.810 2.125 244.240 ;
        RECT 300.170 241.795 301.300 244.225 ;
        RECT 0.995 235.750 2.125 238.180 ;
        RECT 300.170 235.735 301.300 238.165 ;
        RECT 0.995 229.690 2.125 232.120 ;
        RECT 300.170 229.675 301.300 232.105 ;
        RECT 0.995 223.630 2.125 226.060 ;
        RECT 300.170 223.615 301.300 226.045 ;
        RECT 0.995 217.570 2.125 220.000 ;
        RECT 300.170 217.555 301.300 219.985 ;
        RECT 0.995 211.510 2.125 213.940 ;
        RECT 300.170 211.495 301.300 213.925 ;
        RECT 0.995 205.450 2.125 207.880 ;
        RECT 300.170 205.435 301.300 207.865 ;
        RECT 0.995 199.390 2.125 201.820 ;
        RECT 300.170 199.375 301.300 201.805 ;
        RECT 0.995 193.330 2.125 195.760 ;
        RECT 300.170 193.315 301.300 195.745 ;
        RECT 0.995 187.270 2.125 189.700 ;
        RECT 300.170 187.255 301.300 189.685 ;
        RECT 0.995 181.210 2.125 183.640 ;
        RECT 300.170 181.195 301.300 183.625 ;
        RECT 0.995 175.150 2.125 177.580 ;
        RECT 300.170 175.135 301.300 177.565 ;
        RECT 0.995 169.090 2.125 171.520 ;
        RECT 300.170 169.075 301.300 171.505 ;
        RECT 0.995 163.030 2.125 165.460 ;
        RECT 300.170 163.015 301.300 165.445 ;
        RECT 0.995 156.970 2.125 159.400 ;
        RECT 300.170 156.955 301.300 159.385 ;
        RECT 0.995 150.910 2.125 153.340 ;
        RECT 300.170 150.895 301.300 153.325 ;
        RECT 0.995 144.850 2.125 147.280 ;
        RECT 300.170 144.835 301.300 147.265 ;
        RECT 0.995 138.790 2.125 141.220 ;
        RECT 300.170 138.775 301.300 141.205 ;
        RECT 0.995 132.730 2.125 135.160 ;
        RECT 300.170 132.715 301.300 135.145 ;
        RECT 0.995 126.670 2.125 129.100 ;
        RECT 300.170 126.655 301.300 129.085 ;
        RECT 0.995 119.315 2.125 121.745 ;
        RECT 299.185 119.315 300.315 121.745 ;
        RECT 0.995 91.275 2.125 100.865 ;
        RECT 299.185 91.275 300.315 100.865 ;
        RECT 0.995 74.080 2.125 78.180 ;
        RECT 299.185 74.080 300.315 78.180 ;
        RECT 0.995 50.430 2.125 61.980 ;
        RECT 299.185 50.430 300.315 61.980 ;
        RECT 0.995 35.835 2.125 40.005 ;
        RECT 299.185 35.835 300.315 40.005 ;
        RECT 0.995 20.240 2.125 26.580 ;
        RECT 299.185 20.240 300.315 26.580 ;
        RECT 0.995 8.885 2.125 13.055 ;
        RECT 299.185 8.885 300.315 13.055 ;
        RECT 16.245 0.985 19.745 4.485 ;
        RECT 25.040 0.985 25.820 6.000 ;
        RECT 28.600 0.985 29.385 6.000 ;
        RECT 33.045 0.985 36.545 4.485 ;
        RECT 54.045 0.985 57.545 4.485 ;
        RECT 63.850 0.985 64.630 6.000 ;
        RECT 67.410 0.985 68.195 6.000 ;
        RECT 70.845 0.985 74.345 4.485 ;
        RECT 87.000 0.985 87.775 6.000 ;
        RECT 90.555 0.985 91.335 6.000 ;
        RECT 109.630 0.985 113.130 4.485 ;
        RECT 115.575 0.985 119.075 4.485 ;
        RECT 121.905 0.985 125.405 4.485 ;
        RECT 129.495 4.310 130.275 6.000 ;
        RECT 133.055 4.485 133.840 6.000 ;
        RECT 135.865 4.485 136.645 6.000 ;
        RECT 133.055 4.310 136.645 4.485 ;
        RECT 139.425 4.310 140.210 6.000 ;
        RECT 133.095 0.985 136.595 4.310 ;
        RECT 144.315 0.985 147.815 4.485 ;
        RECT 152.715 0.985 156.215 4.485 ;
        RECT 161.115 0.985 164.615 4.485 ;
        RECT 179.315 0.985 182.815 4.485 ;
        RECT 183.670 0.985 187.170 4.485 ;
        RECT 206.100 0.985 206.875 6.000 ;
        RECT 209.655 0.985 210.435 6.000 ;
        RECT 223.760 0.985 227.260 4.485 ;
        RECT 230.315 0.985 231.095 6.000 ;
        RECT 233.875 0.985 234.660 6.000 ;
        RECT 240.560 0.985 244.060 4.485 ;
        RECT 261.560 0.985 265.060 4.485 ;
        RECT 269.465 0.985 270.245 6.000 ;
        RECT 273.025 0.985 273.810 6.000 ;
        RECT 278.360 0.985 281.860 4.485 ;
      LAYER Metal3 ;
        RECT 9.340 327.575 12.840 329.710 ;
        RECT 18.760 327.580 22.265 329.710 ;
        RECT 28.890 327.575 32.390 329.710 ;
        RECT 37.660 327.580 41.165 329.710 ;
        RECT 48.440 327.575 51.940 329.710 ;
        RECT 56.560 327.580 60.065 329.710 ;
        RECT 67.990 327.575 71.490 329.710 ;
        RECT 80.450 329.705 83.950 329.710 ;
        RECT 80.450 327.580 83.960 329.705 ;
        RECT 88.800 327.580 92.305 329.710 ;
        RECT 98.315 327.580 101.820 329.710 ;
        RECT 103.205 327.580 106.705 329.710 ;
        RECT 114.080 327.580 117.585 329.710 ;
        RECT 119.830 327.580 123.335 329.710 ;
        RECT 130.065 327.580 133.570 329.710 ;
        RECT 140.335 327.580 143.840 329.710 ;
        RECT 149.255 327.580 152.755 329.710 ;
        RECT 153.745 327.580 157.245 329.710 ;
        RECT 166.375 327.580 169.880 329.710 ;
        RECT 177.375 327.580 180.880 329.710 ;
        RECT 196.715 327.580 200.215 329.710 ;
        RECT 205.515 328.095 209.020 329.710 ;
        RECT 205.520 327.580 209.020 328.095 ;
        RECT 80.460 327.575 83.960 327.580 ;
        RECT 214.805 327.575 218.305 329.710 ;
        RECT 226.275 327.580 229.780 329.710 ;
        RECT 234.355 329.705 237.855 329.710 ;
        RECT 234.345 327.580 237.855 329.705 ;
        RECT 245.175 327.580 248.680 329.710 ;
        RECT 234.345 327.575 237.845 327.580 ;
        RECT 253.855 327.575 257.355 329.710 ;
        RECT 264.075 327.580 267.580 329.710 ;
        RECT 273.405 327.575 276.905 329.710 ;
        RECT 285.815 329.705 289.315 329.710 ;
        RECT 285.815 327.580 289.325 329.705 ;
        RECT 285.825 327.575 289.325 327.580 ;
        RECT 0.000 322.330 3.555 323.030 ;
        RECT 297.755 322.910 301.300 323.015 ;
        RECT 297.750 322.515 301.300 322.910 ;
        RECT 0.000 321.280 6.000 322.330 ;
        RECT 295.300 321.465 301.300 322.515 ;
        RECT 0.000 320.580 3.555 321.280 ;
        RECT 297.750 320.465 301.300 321.465 ;
        RECT 0.000 316.270 3.555 316.970 ;
        RECT 297.750 316.455 301.300 316.955 ;
        RECT 0.000 315.220 6.000 316.270 ;
        RECT 295.300 315.405 301.300 316.455 ;
        RECT 0.000 314.520 3.555 315.220 ;
        RECT 297.750 314.505 301.300 315.405 ;
        RECT 0.000 310.210 3.555 310.910 ;
        RECT 297.750 310.395 301.300 310.895 ;
        RECT 0.000 309.160 6.000 310.210 ;
        RECT 295.300 309.345 301.300 310.395 ;
        RECT 0.000 308.460 3.555 309.160 ;
        RECT 297.750 308.445 301.300 309.345 ;
        RECT 0.000 304.150 3.555 304.850 ;
        RECT 297.750 304.335 301.300 304.835 ;
        RECT 0.000 303.100 6.000 304.150 ;
        RECT 295.300 303.285 301.300 304.335 ;
        RECT 0.000 302.400 3.555 303.100 ;
        RECT 297.750 302.385 301.300 303.285 ;
        RECT 0.000 298.090 3.555 298.790 ;
        RECT 297.750 298.275 301.300 298.775 ;
        RECT 0.000 297.040 6.000 298.090 ;
        RECT 295.300 297.225 301.300 298.275 ;
        RECT 0.000 296.340 3.555 297.040 ;
        RECT 297.750 296.325 301.300 297.225 ;
        RECT 0.000 292.030 3.555 292.730 ;
        RECT 297.750 292.215 301.300 292.715 ;
        RECT 0.000 290.980 6.000 292.030 ;
        RECT 295.300 291.165 301.300 292.215 ;
        RECT 0.000 290.280 3.555 290.980 ;
        RECT 297.750 290.265 301.300 291.165 ;
        RECT 0.000 285.970 3.555 286.670 ;
        RECT 297.750 286.155 301.300 286.655 ;
        RECT 0.000 284.920 6.000 285.970 ;
        RECT 295.300 285.105 301.300 286.155 ;
        RECT 0.000 284.220 3.555 284.920 ;
        RECT 297.750 284.205 301.300 285.105 ;
        RECT 0.000 279.910 3.555 280.610 ;
        RECT 297.750 280.095 301.300 280.595 ;
        RECT 0.000 278.860 6.000 279.910 ;
        RECT 295.300 279.045 301.300 280.095 ;
        RECT 0.000 278.160 3.555 278.860 ;
        RECT 297.750 278.145 301.300 279.045 ;
        RECT 0.000 273.850 3.555 274.550 ;
        RECT 297.750 274.035 301.300 274.535 ;
        RECT 0.000 272.800 6.000 273.850 ;
        RECT 295.300 272.985 301.300 274.035 ;
        RECT 0.000 272.100 3.555 272.800 ;
        RECT 297.750 272.085 301.300 272.985 ;
        RECT 0.000 267.790 3.555 268.490 ;
        RECT 297.750 267.975 301.300 268.475 ;
        RECT 0.000 266.740 6.000 267.790 ;
        RECT 295.300 266.925 301.300 267.975 ;
        RECT 0.000 266.040 3.555 266.740 ;
        RECT 297.750 266.025 301.300 266.925 ;
        RECT 0.000 261.730 3.555 262.430 ;
        RECT 297.750 261.915 301.300 262.415 ;
        RECT 0.000 260.680 6.000 261.730 ;
        RECT 295.300 260.865 301.300 261.915 ;
        RECT 0.000 259.980 3.555 260.680 ;
        RECT 297.750 259.965 301.300 260.865 ;
        RECT 0.000 255.670 3.555 256.370 ;
        RECT 297.750 255.855 301.300 256.355 ;
        RECT 0.000 254.620 6.000 255.670 ;
        RECT 295.300 254.805 301.300 255.855 ;
        RECT 0.000 253.920 3.555 254.620 ;
        RECT 297.750 253.905 301.300 254.805 ;
        RECT 0.000 249.610 3.555 250.310 ;
        RECT 297.750 249.795 301.300 250.295 ;
        RECT 0.000 248.560 6.000 249.610 ;
        RECT 295.300 248.745 301.300 249.795 ;
        RECT 0.000 247.860 3.555 248.560 ;
        RECT 297.750 247.845 301.300 248.745 ;
        RECT 0.000 243.550 3.555 244.250 ;
        RECT 297.750 243.735 301.300 244.235 ;
        RECT 0.000 242.500 6.000 243.550 ;
        RECT 295.300 242.685 301.300 243.735 ;
        RECT 0.000 241.800 3.555 242.500 ;
        RECT 297.750 241.785 301.300 242.685 ;
        RECT 0.000 237.490 3.555 238.190 ;
        RECT 297.750 237.675 301.300 238.175 ;
        RECT 0.000 236.440 6.000 237.490 ;
        RECT 295.300 236.625 301.300 237.675 ;
        RECT 0.000 235.740 3.555 236.440 ;
        RECT 297.750 235.725 301.300 236.625 ;
        RECT 0.000 231.430 3.555 232.130 ;
        RECT 297.750 231.615 301.300 232.115 ;
        RECT 0.000 230.380 6.000 231.430 ;
        RECT 295.300 230.565 301.300 231.615 ;
        RECT 0.000 229.680 3.555 230.380 ;
        RECT 297.750 229.665 301.300 230.565 ;
        RECT 0.000 225.370 3.555 226.070 ;
        RECT 297.750 225.555 301.300 226.055 ;
        RECT 0.000 224.320 6.000 225.370 ;
        RECT 295.300 224.505 301.300 225.555 ;
        RECT 0.000 223.620 3.555 224.320 ;
        RECT 297.750 223.605 301.300 224.505 ;
        RECT 0.000 219.310 3.555 220.010 ;
        RECT 297.750 219.495 301.300 219.995 ;
        RECT 0.000 218.260 6.000 219.310 ;
        RECT 295.300 218.445 301.300 219.495 ;
        RECT 0.000 217.560 3.555 218.260 ;
        RECT 297.750 217.545 301.300 218.445 ;
        RECT 0.000 213.250 3.555 213.950 ;
        RECT 297.750 213.435 301.300 213.935 ;
        RECT 0.000 212.200 6.000 213.250 ;
        RECT 295.300 212.385 301.300 213.435 ;
        RECT 0.000 211.500 3.555 212.200 ;
        RECT 297.750 211.485 301.300 212.385 ;
        RECT 0.000 207.190 3.555 207.890 ;
        RECT 297.750 207.375 301.300 207.875 ;
        RECT 0.000 206.140 6.000 207.190 ;
        RECT 295.300 206.325 301.300 207.375 ;
        RECT 0.000 205.440 3.555 206.140 ;
        RECT 297.750 205.425 301.300 206.325 ;
        RECT 0.000 201.130 3.555 201.830 ;
        RECT 297.750 201.315 301.300 201.815 ;
        RECT 0.000 200.080 6.000 201.130 ;
        RECT 295.300 200.265 301.300 201.315 ;
        RECT 0.000 199.380 3.555 200.080 ;
        RECT 297.750 199.365 301.300 200.265 ;
        RECT 0.000 195.070 3.555 195.770 ;
        RECT 297.750 195.255 301.300 195.755 ;
        RECT 0.000 194.020 6.000 195.070 ;
        RECT 295.300 194.205 301.300 195.255 ;
        RECT 0.000 193.320 3.555 194.020 ;
        RECT 297.750 193.305 301.300 194.205 ;
        RECT 0.000 189.010 3.555 189.710 ;
        RECT 297.750 189.195 301.300 189.695 ;
        RECT 0.000 187.960 6.000 189.010 ;
        RECT 295.300 188.145 301.300 189.195 ;
        RECT 0.000 187.260 3.555 187.960 ;
        RECT 297.750 187.245 301.300 188.145 ;
        RECT 0.000 182.950 3.555 183.650 ;
        RECT 297.750 183.135 301.300 183.635 ;
        RECT 0.000 181.900 6.000 182.950 ;
        RECT 295.300 182.085 301.300 183.135 ;
        RECT 0.000 181.200 3.555 181.900 ;
        RECT 297.750 181.185 301.300 182.085 ;
        RECT 0.000 176.890 3.555 177.590 ;
        RECT 297.750 177.075 301.300 177.575 ;
        RECT 0.000 175.840 6.000 176.890 ;
        RECT 295.300 176.025 301.300 177.075 ;
        RECT 0.000 175.140 3.555 175.840 ;
        RECT 297.750 175.125 301.300 176.025 ;
        RECT 0.000 170.830 3.555 171.530 ;
        RECT 297.750 171.015 301.300 171.515 ;
        RECT 0.000 169.780 6.000 170.830 ;
        RECT 295.300 169.965 301.300 171.015 ;
        RECT 0.000 169.080 3.555 169.780 ;
        RECT 297.750 169.065 301.300 169.965 ;
        RECT 0.000 164.770 3.555 165.470 ;
        RECT 297.750 164.955 301.300 165.455 ;
        RECT 0.000 163.720 6.000 164.770 ;
        RECT 295.300 163.905 301.300 164.955 ;
        RECT 0.000 163.020 3.555 163.720 ;
        RECT 297.750 163.005 301.300 163.905 ;
        RECT 0.000 158.710 3.555 159.410 ;
        RECT 297.750 158.895 301.300 159.395 ;
        RECT 0.000 157.660 6.000 158.710 ;
        RECT 295.300 157.845 301.300 158.895 ;
        RECT 0.000 156.960 3.555 157.660 ;
        RECT 297.750 156.945 301.300 157.845 ;
        RECT 0.000 152.650 3.555 153.350 ;
        RECT 297.750 152.835 301.300 153.335 ;
        RECT 0.000 151.600 6.000 152.650 ;
        RECT 295.300 151.785 301.300 152.835 ;
        RECT 0.000 150.900 3.555 151.600 ;
        RECT 297.750 150.885 301.300 151.785 ;
        RECT 0.000 146.590 3.555 147.290 ;
        RECT 297.750 146.775 301.300 147.275 ;
        RECT 0.000 145.540 6.000 146.590 ;
        RECT 295.300 145.725 301.300 146.775 ;
        RECT 0.000 144.840 3.555 145.540 ;
        RECT 297.750 144.825 301.300 145.725 ;
        RECT 0.000 140.530 3.555 141.230 ;
        RECT 297.750 140.715 301.300 141.215 ;
        RECT 0.000 139.480 6.000 140.530 ;
        RECT 295.300 139.665 301.300 140.715 ;
        RECT 0.000 138.780 3.555 139.480 ;
        RECT 297.750 138.765 301.300 139.665 ;
        RECT 0.000 134.470 3.555 135.170 ;
        RECT 297.755 135.010 301.300 135.155 ;
        RECT 297.750 134.655 301.300 135.010 ;
        RECT 0.000 133.420 6.000 134.470 ;
        RECT 295.300 133.605 301.300 134.655 ;
        RECT 0.000 132.720 3.555 133.420 ;
        RECT 297.750 132.705 301.300 133.605 ;
        RECT 0.000 128.410 3.555 129.110 ;
        RECT 297.755 128.900 301.300 129.095 ;
        RECT 297.750 128.595 301.300 128.900 ;
        RECT 0.000 127.360 6.000 128.410 ;
        RECT 295.300 127.545 301.300 128.595 ;
        RECT 0.000 126.660 3.555 127.360 ;
        RECT 297.750 126.645 301.300 127.545 ;
        RECT 0.010 121.935 6.000 122.180 ;
        RECT 0.000 121.480 6.000 121.935 ;
        RECT 295.300 121.480 301.300 122.180 ;
        RECT 0.000 120.845 3.555 121.480 ;
        RECT 297.750 120.845 301.300 121.480 ;
        RECT 0.000 119.170 6.000 120.845 ;
        RECT 0.010 119.165 6.000 119.170 ;
        RECT 295.300 119.165 301.300 120.845 ;
        RECT 0.000 100.995 3.545 101.000 ;
        RECT 297.750 100.995 301.300 101.000 ;
        RECT 0.000 94.065 6.000 100.995 ;
        RECT 0.010 94.060 6.000 94.065 ;
        RECT 295.300 94.060 301.300 100.995 ;
        RECT 295.300 94.045 295.500 94.060 ;
        RECT 0.000 78.275 3.545 78.280 ;
        RECT 297.755 78.275 301.300 78.280 ;
        RECT 0.000 76.685 6.000 78.275 ;
        RECT 295.300 76.685 301.300 78.275 ;
        RECT 0.000 74.780 3.555 76.685 ;
        RECT 295.300 76.680 295.315 76.685 ;
        RECT 297.755 76.280 301.300 76.685 ;
        RECT 297.750 74.780 301.300 76.280 ;
        RECT 0.010 74.775 3.555 74.780 ;
        RECT 297.755 74.775 301.300 74.780 ;
        RECT 0.000 62.045 3.545 62.100 ;
        RECT 297.750 62.045 301.300 62.050 ;
        RECT 0.000 50.190 6.000 62.045 ;
        RECT 0.010 50.135 6.000 50.190 ;
        RECT 295.300 50.135 301.300 62.045 ;
        RECT 0.000 40.215 3.545 40.270 ;
        RECT 297.750 40.215 301.300 40.220 ;
        RECT 0.000 35.660 6.000 40.215 ;
        RECT 0.010 35.605 6.000 35.660 ;
        RECT 295.300 35.605 301.300 40.215 ;
        RECT 0.000 26.575 3.545 26.630 ;
        RECT 297.750 26.575 301.300 26.580 ;
        RECT 0.000 24.425 6.000 26.575 ;
        RECT 295.300 24.425 301.300 26.575 ;
        RECT 0.000 21.685 3.555 24.425 ;
        RECT 295.300 24.420 295.750 24.425 ;
        RECT 297.750 21.685 301.300 24.425 ;
        RECT 0.000 20.225 6.000 21.685 ;
        RECT 0.010 20.170 6.000 20.225 ;
        RECT 295.300 20.170 301.300 21.685 ;
        RECT 0.000 13.190 3.545 13.245 ;
        RECT 300.600 13.190 301.300 13.195 ;
        RECT 0.000 11.960 6.000 13.190 ;
        RECT 295.300 11.960 301.300 13.190 ;
        RECT 0.000 10.030 3.545 11.960 ;
        RECT 297.805 11.495 301.300 11.960 ;
        RECT 297.750 10.030 301.300 11.495 ;
        RECT 0.000 8.800 6.000 10.030 ;
        RECT 0.010 8.745 6.000 8.800 ;
        RECT 295.300 8.745 301.300 10.030 ;
        RECT 16.245 0.000 19.745 3.260 ;
        RECT 33.045 0.000 36.545 3.260 ;
        RECT 54.045 0.000 57.545 3.260 ;
        RECT 70.845 0.000 74.345 3.260 ;
        RECT 109.630 0.000 113.130 3.260 ;
        RECT 115.575 0.000 119.075 3.260 ;
        RECT 121.905 0.000 125.405 3.260 ;
        RECT 133.095 0.000 136.595 3.260 ;
        RECT 144.315 0.000 147.815 3.260 ;
        RECT 152.715 0.000 156.215 3.260 ;
        RECT 161.115 0.000 164.615 3.260 ;
        RECT 179.315 0.000 182.815 3.260 ;
        RECT 183.670 0.000 187.170 3.260 ;
        RECT 223.760 0.000 227.260 3.260 ;
        RECT 240.560 0.000 244.060 3.260 ;
        RECT 261.560 0.000 265.060 3.260 ;
        RECT 278.360 0.000 281.860 3.260 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.738400 ;
    PORT
      LAYER Metal2 ;
        RECT 97.775 0.000 98.560 6.000 ;
    END
  END CLK
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 6.520 0.000 7.305 6.000 ;
    END
  END D[0]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 101.520 0.000 102.305 6.000 ;
    END
  END A[8]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 103.965 0.000 104.750 6.000 ;
    END
  END A[7]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 108.005 0.000 108.790 6.000 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 113.930 0.000 114.715 6.000 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 119.850 0.000 120.630 6.000 ;
    END
  END A[0]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 51.250 5.450 51.580 6.000 ;
        RECT 49.960 5.120 51.580 5.450 ;
        RECT 49.960 4.160 50.290 5.120 ;
        RECT 49.440 3.710 50.290 4.160 ;
        RECT 49.440 0.000 50.225 3.710 ;
    END
  END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 77.980 4.130 78.315 6.000 ;
        RECT 77.975 0.000 78.760 4.130 ;
    END
  END Q[3]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 176.195 0.000 176.980 6.000 ;
    END
  END CEN
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 190.455 0.000 191.240 6.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 188.200 0.000 188.985 6.000 ;
    END
  END A[6]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 193.070 0.000 193.855 6.000 ;
    END
  END A[4]
  PIN WEN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 81.990 5.975 82.620 5.990 ;
        RECT 81.990 5.945 84.110 5.975 ;
        RECT 81.990 5.685 84.470 5.945 ;
        RECT 81.990 5.670 84.110 5.685 ;
        RECT 81.990 5.650 82.620 5.670 ;
      LAYER Metal2 ;
        RECT 81.910 0.000 82.695 6.000 ;
    END
  END WEN[3]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 291.200 5.030 291.985 6.000 ;
        RECT 290.800 4.305 291.985 5.030 ;
        RECT 290.800 0.000 291.585 4.305 ;
    END
  END D[7]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 285.870 4.245 286.200 6.000 ;
        RECT 285.490 0.000 286.275 4.245 ;
    END
  END Q[7]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 83.280 4.350 84.065 4.380 ;
        RECT 85.695 4.350 86.000 6.000 ;
        RECT 83.280 4.045 86.000 4.350 ;
        RECT 83.280 0.000 84.065 4.045 ;
    END
  END D[3]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 43.215 4.600 43.540 6.000 ;
        RECT 43.180 4.170 43.540 4.600 ;
        RECT 42.720 0.000 43.505 4.170 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 48.730 5.425 49.015 6.000 ;
        RECT 47.595 5.140 49.015 5.425 ;
        RECT 47.595 4.160 47.880 5.140 ;
        RECT 47.085 3.720 47.880 4.160 ;
        RECT 47.085 0.000 47.870 3.720 ;
    END
  END D[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 196.925 0.000 197.710 6.000 ;
    END
  END A[3]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 41.545 4.725 41.875 6.000 ;
        RECT 40.840 4.395 41.875 4.725 ;
        RECT 40.840 4.200 41.170 4.395 ;
        RECT 40.365 3.555 41.170 4.200 ;
        RECT 40.365 0.000 41.145 3.555 ;
    END
  END Q[1]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 257.025 4.245 257.345 6.000 ;
        RECT 256.960 0.000 257.740 4.245 ;
    END
  END Q[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 249.530 4.245 249.810 6.000 ;
        RECT 249.235 0.000 250.020 4.245 ;
    END
  END D[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 217.860 4.705 218.190 6.000 ;
        RECT 217.860 4.695 220.060 4.705 ;
        RECT 217.860 4.375 220.135 4.695 ;
        RECT 219.350 0.000 220.135 4.375 ;
    END
  END Q[4]
  PIN WEN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 249.780 5.945 250.340 5.975 ;
        RECT 250.710 5.945 251.340 5.985 ;
        RECT 249.775 5.685 251.340 5.945 ;
        RECT 249.780 5.675 250.340 5.685 ;
        RECT 250.710 5.645 251.340 5.685 ;
      LAYER Metal2 ;
        RECT 250.630 0.000 251.410 6.000 ;
    END
  END WEN[5]
  PIN WEN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 45.915 5.940 46.545 5.990 ;
        RECT 48.235 5.945 48.795 5.975 ;
        RECT 47.630 5.940 48.800 5.945 ;
        RECT 45.915 5.685 48.800 5.940 ;
        RECT 45.915 5.675 48.795 5.685 ;
        RECT 45.915 5.665 48.390 5.675 ;
        RECT 45.915 5.650 46.545 5.665 ;
      LAYER Metal2 ;
        RECT 45.685 5.650 46.545 5.990 ;
        RECT 45.685 0.000 46.470 5.650 ;
    END
  END WEN[2]
  PIN WEN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 44.190 5.975 44.820 5.990 ;
        RECT 44.190 5.945 45.035 5.975 ;
        RECT 44.190 5.685 45.640 5.945 ;
        RECT 44.190 5.675 45.035 5.685 ;
        RECT 44.190 5.665 44.945 5.675 ;
        RECT 44.190 5.650 44.820 5.665 ;
      LAYER Metal2 ;
        RECT 44.110 0.000 44.895 5.995 ;
    END
  END WEN[1]
  PIN WEN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 214.710 5.950 215.270 5.975 ;
        RECT 214.320 5.945 216.880 5.950 ;
        RECT 214.105 5.940 216.880 5.945 ;
        RECT 214.105 5.690 217.110 5.940 ;
        RECT 214.105 5.685 215.275 5.690 ;
        RECT 214.710 5.675 215.270 5.685 ;
        RECT 216.480 5.600 217.110 5.690 ;
      LAYER Metal2 ;
        RECT 216.400 0.000 217.185 5.955 ;
    END
  END WEN[4]
  PIN WEN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 288.510 5.980 289.140 5.990 ;
        RECT 288.510 5.950 289.420 5.980 ;
        RECT 288.510 5.690 290.025 5.950 ;
        RECT 288.510 5.680 289.420 5.690 ;
        RECT 288.510 5.650 289.140 5.680 ;
      LAYER Metal2 ;
        RECT 288.430 0.000 289.215 5.995 ;
    END
  END WEN[7]
  PIN WEN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 253.285 5.980 253.915 5.985 ;
        RECT 253.285 5.950 254.350 5.980 ;
        RECT 253.185 5.690 254.355 5.950 ;
        RECT 253.285 5.680 254.350 5.690 ;
        RECT 253.285 5.645 253.915 5.680 ;
      LAYER Metal2 ;
        RECT 253.205 0.000 253.985 6.000 ;
    END
  END WEN[6]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 212.255 4.355 212.625 6.000 ;
        RECT 212.255 3.985 214.845 4.355 ;
        RECT 214.060 0.000 214.845 3.985 ;
    END
  END D[4]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 254.645 4.245 254.930 6.000 ;
        RECT 254.605 0.000 255.385 4.245 ;
    END
  END D[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 247.175 4.245 247.460 6.000 ;
        RECT 246.880 0.000 247.665 4.245 ;
    END
  END Q[5]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 12.255 4.245 12.585 6.000 ;
        RECT 11.830 0.000 12.610 4.245 ;
    END
  END Q[0]
  PIN GWEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.141600 ;
    PORT
      LAYER Metal2 ;
        RECT 142.055 0.000 142.840 6.000 ;
    END
  END GWEN
  PIN WEN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.965 5.975 9.595 5.985 ;
        RECT 8.965 5.945 9.965 5.975 ;
        RECT 8.800 5.685 9.970 5.945 ;
        RECT 8.965 5.675 9.965 5.685 ;
        RECT 8.965 5.645 9.595 5.675 ;
      LAYER Metal2 ;
        RECT 8.965 5.980 9.595 5.985 ;
        RECT 8.885 0.000 9.670 5.980 ;
    END
  END WEN[0]
  OBS
      LAYER Nwell ;
        RECT 6.305 6.000 295.010 323.865 ;
      LAYER Metal1 ;
        RECT 6.000 6.000 295.300 323.865 ;
      LAYER Metal2 ;
        RECT 6.000 6.000 295.300 323.865 ;
      LAYER Metal3 ;
        RECT 6.000 93.570 295.300 323.865 ;
        RECT 6.000 92.820 295.500 93.570 ;
        RECT 6.000 92.345 295.300 92.820 ;
        RECT 6.000 91.590 295.500 92.345 ;
        RECT 6.000 91.120 295.300 91.590 ;
        RECT 6.000 90.365 295.500 91.120 ;
        RECT 6.000 89.895 295.300 90.365 ;
        RECT 6.000 89.140 295.500 89.895 ;
        RECT 6.000 6.000 295.300 89.140 ;
  END
END gf180mcu_ocd_ip_sram__sram512x8m8wm1
END LIBRARY

