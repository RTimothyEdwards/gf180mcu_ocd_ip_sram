magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal1 >>
rect 103 52 218 1209
<< metal2 >>
rect 252 0 322 983
<< metal3 >>
rect -357 437 342 1697
rect 499 1271 1199 1697
use M2_M14310591302017_256x8m81  M2_M14310591302017_256x8m81_0
timestamp 1763766357
transform 1 0 849 0 1 1386
box -330 -113 330 113
use M3_M24310591302016_256x8m81  M3_M24310591302016_256x8m81_0
timestamp 1763766357
transform 1 0 849 0 1 1386
box -330 -113 330 113
use M3_M24310591302042_256x8m81  M3_M24310591302042_256x8m81_0
timestamp 1763766357
transform 1 0 -8 0 1 788
box -330 -330 330 330
<< properties >>
string path -0.055 12.125 -0.055 3.125 
<< end >>
