magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< error_s >>
rect 15338 2703 15349 2706
rect 15394 2341 15405 2703
rect 623 1808 662 1809
rect 696 1808 735 1809
rect 821 1808 860 1809
rect 894 1808 933 1809
rect 1019 1808 1058 1809
rect 1092 1808 1131 1809
rect 1903 1808 1942 1809
rect 1976 1808 2015 1809
rect 2101 1808 2140 1809
rect 2174 1808 2213 1809
rect 2299 1808 2338 1809
rect 2372 1808 2411 1809
rect 5788 1808 5827 1809
rect 5861 1808 5900 1809
rect 5986 1808 6025 1809
rect 6059 1808 6098 1809
rect 6184 1808 6223 1809
rect 6257 1808 6296 1809
rect 7068 1808 7107 1809
rect 7141 1808 7180 1809
rect 7266 1808 7305 1809
rect 7339 1808 7378 1809
rect 7464 1808 7503 1809
rect 7537 1808 7576 1809
<< nwell >>
rect 5166 5590 5233 5782
rect 5166 5302 5374 5590
rect 5170 3963 5374 5302
<< metal2 >>
rect 684 7739 775 7833
rect 933 7739 1024 7833
rect 1937 7739 2028 7833
rect 2191 7739 2282 7833
rect 2875 7135 3123 8738
rect 3650 7340 3740 8019
rect 5849 7739 5940 7833
rect 6099 7739 6189 7833
rect 7102 7739 7193 7833
rect 7356 7739 7446 7833
rect 8815 7340 8905 8019
rect 10497 8005 10744 8780
rect 9007 7750 10744 8005
rect 9007 7134 9254 7750
rect 11028 7506 11183 7991
rect 11274 7506 11429 7991
rect 12172 7506 12327 7991
rect 12418 7506 12573 7991
rect 13316 7506 13471 7991
rect 13561 7506 13717 7991
rect 14459 7506 14614 7991
rect 14705 7506 14861 7991
rect 15210 7508 15457 8738
rect 16135 7604 16226 8019
rect 15210 7415 15544 7508
rect 15422 7414 15544 7415
rect 16344 2048 16434 2142
rect 17528 2048 17618 2142
rect 18711 2048 18802 2142
rect 3857 1854 3947 1948
rect 5041 1854 5131 1948
rect 9022 1854 9113 1948
rect 10205 1854 10296 1948
<< metal3 >>
rect 32 8145 19082 8780
rect 32 7843 15349 8060
rect 5256 2787 5777 3265
rect 5256 2340 5777 2705
rect 5256 1813 5777 2267
use M3_M2$$43368492_3v512x8m81  M3_M2$$43368492_3v512x8m81_0
timestamp 1763765945
transform 1 0 3695 0 1 7966
box -44 -123 44 123
use M3_M2$$43368492_3v512x8m81  M3_M2$$43368492_3v512x8m81_1
timestamp 1763765945
transform 0 1 8783 -1 0 7976
box -44 -123 44 123
use M3_M2$$43368492_3v512x8m81  M3_M2$$43368492_3v512x8m81_2
timestamp 1763765945
transform 0 1 16259 -1 0 7971
box -44 -123 44 123
use M3_M2$$47115308_3v512x8m81  M3_M2$$47115308_3v512x8m81_0
timestamp 1763765945
transform 1 0 2979 0 1 8463
box -119 -275 119 275
use M3_M2$$47115308_3v512x8m81  M3_M2$$47115308_3v512x8m81_1
timestamp 1763765945
transform 1 0 15334 0 1 8463
box -119 -275 119 275
use M3_M2$$201412652_3v512x8m81  M3_M2$$201412652_3v512x8m81_0
timestamp 1763765945
transform 1 0 10620 0 1 8463
box -119 -275 119 275
use xpredec0_3v512x8m81  xpredec0_3v512x8m81_0
timestamp 1763765945
transform 1 0 5412 0 1 0
box -226 1806 10233 8019
use xpredec0_3v512x8m81  xpredec0_3v512x8m81_1
timestamp 1763765945
transform 1 0 247 0 1 0
box -226 1806 10233 8019
use xpredec1_3v512x8m81  xpredec1_3v512x8m81_0
timestamp 1763765945
transform 1 0 10557 0 1 400
box -1 1414 8563 7679
<< labels >>
rlabel metal3 s 17852 8463 17852 8463 4 men
port 2 nsew
rlabel metal2 s 5895 7786 5895 7786 4 xb[3]
port 6 nsew
rlabel metal2 s 14786 7945 14786 7945 4 xa[0]
port 7 nsew
rlabel metal2 s 2236 7784 2236 7784 4 xc[0]
port 8 nsew
rlabel metal2 s 1983 7784 1983 7784 4 xc[1]
port 9 nsew
rlabel metal2 s 979 7786 979 7786 4 xc[2]
port 10 nsew
rlabel metal2 s 730 7786 730 7786 4 xc[3]
port 11 nsew
rlabel metal2 s 7147 7784 7147 7784 4 xb[1]
port 12 nsew
rlabel metal2 s 6143 7786 6143 7786 4 xb[2]
port 13 nsew
rlabel metal2 s 7401 7784 7401 7784 4 xb[0]
port 14 nsew
rlabel metal2 s 14534 7945 14534 7945 4 xa[1]
port 15 nsew
rlabel metal2 s 13633 7945 13633 7945 4 xa[2]
port 16 nsew
rlabel metal2 s 13393 7945 13393 7945 4 xa[3]
port 17 nsew
rlabel metal2 s 12497 7945 12497 7945 4 xa[4]
port 18 nsew
rlabel metal2 s 12248 7945 12248 7945 4 xa[5]
port 19 nsew
rlabel metal2 s 11350 7945 11350 7945 4 xa[6]
port 20 nsew
rlabel metal2 s 11104 7945 11104 7945 4 xa[7]
port 21 nsew
rlabel metal2 s 3902 1901 3902 1901 4 A[6]
port 4 nsew
rlabel metal2 s 9067 1901 9067 1901 4 A[4]
port 5 nsew
rlabel metal2 s 10251 1901 10251 1901 4 A[3]
port 23 nsew
rlabel metal2 s 5086 1901 5086 1901 4 A[5]
port 24 nsew
rlabel metal2 s 16389 2095 16389 2095 4 A[2]
port 3 nsew
rlabel metal2 s 17573 2095 17573 2095 4 A[1]
port 25 nsew
rlabel metal2 s 18757 2095 18757 2095 4 A[0]
port 22 nsew
<< end >>
