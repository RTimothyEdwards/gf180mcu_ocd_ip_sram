magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal2 >>
rect -330 323 330 330
rect -330 -323 -323 323
rect 323 -323 330 323
rect -330 -330 330 -323
<< via2 >>
rect -323 -323 323 323
<< metal3 >>
rect -330 323 330 330
rect -330 -323 -323 323
rect 323 -323 330 323
rect -330 -330 330 -323
<< end >>
