magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_0
timestamp 1763564386
transform 1 0 0 0 1 0
box -8 0 72 215
use via2_x2_R90_512x8m81  via2_x2_R90_512x8m81_0
timestamp 1763564386
transform 1 0 0 0 1 0
box -9 0 73 215
<< end >>
