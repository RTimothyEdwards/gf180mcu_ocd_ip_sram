magic
tech gf180mcuD
magscale 1 10
timestamp 1763255117
<< metal1 >>
rect -44 26 45 46
rect -44 -26 -26 26
rect 26 -26 45 26
rect -44 -46 45 -26
<< via1 >>
rect -26 -26 26 26
<< metal2 >>
rect -44 26 45 46
rect -44 -26 -26 26
rect 26 -26 45 26
rect -44 -46 45 -26
<< end >>
