magic
tech gf180mcuD
magscale 1 10
timestamp 1764092614
<< metal2 >>
rect 1304 0 1461 140
rect 2017 0 2174 140
rect 2766 0 2922 140
rect 8073 0 8229 140
rect 8544 0 8701 140
rect 8822 0 8979 140
rect 9137 0 9294 140
rect 9417 0 9574 140
rect 9888 0 10045 140
rect 15595 0 15752 140
rect 16382 0 16539 140
rect 16656 0 16813 140
rect 19555 0 19712 140
rect 20792 0 20949 140
rect 21601 0 21758 140
rect 22786 0 22943 140
rect 23970 0 24126 140
rect 28411 0 28568 140
rect 35239 0 35396 140
rect 37640 0 37797 140
rect 38091 0 38248 140
rect 38614 0 38771 140
rect 39385 0 39542 140
rect 42812 0 42969 140
rect 43280 0 43437 140
rect 43870 0 44027 140
rect 49376 0 49533 140
rect 49847 0 50004 140
rect 50126 0 50282 140
rect 50641 0 50797 140
rect 50921 0 51077 140
rect 51392 0 51548 140
rect 57098 0 57255 140
rect 57686 0 57843 140
rect 58160 0 58317 140
<< metal3 >>
rect 1010 44846 1710 44986
rect 1868 44846 2568 44986
rect 2895 44846 3595 44986
rect 3753 44846 4453 44986
rect 4920 44846 5620 44986
rect 5778 44846 6478 44986
rect 6675 44846 7375 44986
rect 7533 44846 8233 44986
rect 8830 44846 9530 44986
rect 9688 44846 10388 44986
rect 10455 44846 11155 44986
rect 11313 44846 12013 44986
rect 12740 44846 13440 44986
rect 13598 44846 14298 44986
rect 14457 44846 15157 44986
rect 16090 44846 16790 44986
rect 16948 44846 17648 44986
rect 17760 44846 18460 44986
rect 18600 44846 19300 44986
rect 19663 44846 20363 44986
rect 20641 44846 21341 44986
rect 21497 44846 22197 44986
rect 22816 44846 23516 44986
rect 23966 44846 24666 44986
rect 24790 44846 25490 44986
rect 26013 44846 26713 44986
rect 27009 44846 27709 44986
rect 28067 44846 28767 44986
rect 28861 44846 29561 44986
rect 29851 44846 30551 44986
rect 30749 44846 31449 44986
rect 31548 44846 32248 44986
rect 32419 44846 33119 44986
rect 33276 44846 33976 44986
rect 34230 44846 34930 44986
rect 35475 44846 36175 44986
rect 36798 44846 37498 44986
rect 37983 44846 38683 44986
rect 39343 44846 40043 44986
rect 40282 44846 40982 44986
rect 41103 44846 41803 44986
rect 42103 44846 42803 44986
rect 42961 44846 43661 44986
rect 44399 44846 45099 44986
rect 45256 44846 45956 44986
rect 46013 44846 46713 44986
rect 46871 44846 47571 44986
rect 48179 44846 48879 44986
rect 49036 44846 49736 44986
rect 49913 44846 50613 44986
rect 50771 44846 51471 44986
rect 51959 44846 52659 44986
rect 52816 44846 53516 44986
rect 53823 44846 54523 44986
rect 54681 44846 55381 44986
rect 55860 44846 56560 44986
rect 57163 44846 57863 44986
rect 58021 44846 58721 44986
rect 59066 44846 59766 44986
rect 0 43742 140 44232
rect 60120 43759 60260 44249
rect 0 43160 140 43650
rect 60120 43157 60260 43647
rect 0 42530 140 43020
rect 60120 42547 60260 43037
rect 0 41948 140 42438
rect 60120 41945 60260 42435
rect 0 41318 140 41808
rect 60120 41335 60260 41825
rect 0 40736 140 41226
rect 60120 40733 60260 41223
rect 0 40106 140 40596
rect 60120 40123 60260 40613
rect 0 39524 140 40014
rect 60120 39521 60260 40011
rect 0 38894 140 39384
rect 60120 38911 60260 39401
rect 0 38312 140 38802
rect 60120 38309 60260 38799
rect 0 37682 140 38172
rect 60120 37699 60260 38189
rect 0 37100 140 37590
rect 60120 37097 60260 37587
rect 0 36470 140 36960
rect 60120 36487 60260 36977
rect 0 35888 140 36378
rect 60120 35885 60260 36375
rect 0 35258 140 35748
rect 60120 35275 60260 35765
rect 0 34676 140 35166
rect 60120 34673 60260 35163
rect 0 34046 140 34536
rect 60120 34063 60260 34553
rect 0 33464 140 33954
rect 60120 33461 60260 33951
rect 0 32834 140 33324
rect 60120 32851 60260 33341
rect 0 32252 140 32742
rect 60120 32249 60260 32739
rect 0 31622 140 32112
rect 60120 31639 60260 32129
rect 0 31040 140 31530
rect 60120 31037 60260 31527
rect 0 30410 140 30900
rect 60120 30427 60260 30917
rect 0 29828 140 30318
rect 60120 29825 60260 30315
rect 0 29198 140 29688
rect 60120 29215 60260 29705
rect 0 28616 140 29106
rect 60120 28613 60260 29103
rect 0 27986 140 28476
rect 60120 28003 60260 28493
rect 0 27404 140 27894
rect 60120 27401 60260 27891
rect 0 26774 140 27264
rect 60120 26791 60260 27281
rect 0 26192 140 26682
rect 60120 26189 60260 26679
rect 0 25562 140 26052
rect 60120 25579 60260 26069
rect 0 24980 140 25470
rect 60120 24977 60260 25467
rect 0 24350 140 24840
rect 60120 24367 60260 24857
rect 0 23768 140 24258
rect 60120 23765 60260 24255
rect 0 23138 140 23628
rect 60120 23155 60260 23645
rect 0 22270 140 22823
rect 60120 22270 60260 22823
rect 0 19035 140 21982
rect 60120 19034 60260 21982
rect 0 17379 140 18766
rect 60120 17379 60260 18766
rect 0 14971 140 15671
rect 60120 14971 60260 15671
rect 0 13872 140 14572
rect 60120 13872 60260 14572
rect 0 11641 140 13547
rect 60120 11641 60260 13547
rect 0 9594 140 11441
rect 60120 9590 60260 11441
rect 0 8026 140 9464
rect 60120 8003 60260 9464
rect 0 6723 140 7645
rect 60120 6723 60260 7645
rect 0 5306 140 6260
rect 60120 5306 60260 6260
rect 0 3962 140 5092
rect 60120 3962 60260 5092
rect 0 2842 140 3870
rect 60120 2841 60260 3870
rect 0 1751 140 2640
rect 60120 1750 60260 2639
rect 0 858 140 1558
rect 60120 862 60260 1562
rect 494 0 1194 140
rect 1427 0 2127 140
rect 2409 0 3109 140
rect 3249 0 3949 140
rect 4089 0 4789 140
rect 4929 0 5629 140
rect 5769 0 6469 140
rect 6609 0 7309 140
rect 7449 0 8149 140
rect 8710 0 9410 140
rect 9969 0 10669 140
rect 10809 0 11509 140
rect 11649 0 12349 140
rect 12489 0 13189 140
rect 13329 0 14029 140
rect 14169 0 14869 140
rect 15337 0 16037 140
rect 16177 0 16877 140
rect 17087 0 17787 140
rect 17997 0 18697 140
rect 18907 0 19607 140
rect 19817 0 20517 140
rect 20727 0 21427 140
rect 21926 0 22626 140
rect 23115 0 23815 140
rect 24381 0 25081 140
rect 25221 0 25921 140
rect 26619 0 27319 140
rect 27459 0 28159 140
rect 28863 0 29563 140
rect 29703 0 30403 140
rect 30543 0 31243 140
rect 31383 0 32083 140
rect 32223 0 32923 140
rect 33063 0 33763 140
rect 33996 0 34696 140
rect 34913 0 35613 140
rect 35863 0 36563 140
rect 36734 0 37434 140
rect 38120 0 38820 140
rect 39030 0 39730 140
rect 39940 0 40640 140
rect 40850 0 41550 140
rect 41760 0 42460 140
rect 42670 0 43370 140
rect 43606 0 44306 140
rect 44752 0 45452 140
rect 45592 0 46292 140
rect 46432 0 47132 140
rect 47272 0 47972 140
rect 48112 0 48812 140
rect 48952 0 49652 140
rect 50211 0 50911 140
rect 51472 0 52172 140
rect 52312 0 53012 140
rect 53152 0 53852 140
rect 53992 0 54692 140
rect 54832 0 55532 140
rect 55672 0 56372 140
rect 56712 0 57412 140
rect 57693 0 58393 140
rect 59066 0 59766 140
<< labels >>
flabel metal3 s 70 24058 70 24058 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 23383 70 23383 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 22520 70 22520 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 20858 70 20858 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 24595 70 24595 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 25807 70 25807 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 27019 70 27019 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 28231 70 28231 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 29443 70 29443 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 30655 70 30655 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 31867 70 31867 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 33079 70 33079 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 34291 70 34291 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 35503 70 35503 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 36715 70 36715 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 37927 70 37927 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 39139 70 39139 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 40351 70 40351 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 41563 70 41563 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 42775 70 42775 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 43987 70 43987 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 25222 70 25222 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 26434 70 26434 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 27646 70 27646 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 28858 70 28858 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 30070 70 30070 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 31282 70 31282 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 32494 70 32494 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 33706 70 33706 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 34918 70 34918 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 36130 70 36130 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 37342 70 37342 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 38554 70 38554 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 39766 70 39766 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 40978 70 40978 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 42190 70 42190 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 43402 70 43402 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 22520 60196 22520 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 20858 60196 20858 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 25267 60196 25267 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 24055 60196 24055 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 26479 60196 26479 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 27691 60196 27691 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 28903 60196 28903 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 30115 60196 30115 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 31327 60196 31327 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 32539 60196 32539 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 33751 60196 33751 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 34963 60196 34963 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 36175 60196 36175 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 37387 60196 37387 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 38599 60196 38599 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 39811 60196 39811 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 41023 60196 41023 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 42235 60196 42235 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 43447 60196 43447 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 44004 60196 44004 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 42792 60196 42792 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 41580 60196 41580 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 40368 60196 40368 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 39156 60196 39156 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 37944 60196 37944 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 36732 60196 36732 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 35520 60196 35520 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 34308 60196 34308 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 33096 60196 33096 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 31884 60196 31884 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 30672 60196 30672 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 29460 60196 29460 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 28248 60196 28248 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 27036 60196 27036 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 25824 60196 25824 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 24612 60196 24612 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 23400 60196 23400 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 18236 70 18236 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 15311 70 15311 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 14401 70 14401 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 10254 70 10254 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 11783 70 11783 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 8107 70 8107 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 5448 70 5448 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 7039 70 7039 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 4392 70 4392 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 2914 70 2914 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 70 2214 70 2214 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 70 1178 70 1178 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 18236 60196 18236 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 15311 60196 15311 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 14401 60196 14401 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 10254 60196 10254 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 11783 60196 11783 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 8107 60196 8107 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 7039 60196 7039 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 5757 60196 5757 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 4392 60196 4392 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 3320 60196 3320 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 60196 2213 60196 2213 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 60196 1182 60196 1182 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 2759 70 2759 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 22276 70 22276 70 0 FreeSans 280 180 0 0 VSS
port 1 nsew
flabel metal3 s 23464 70 23464 70 0 FreeSans 280 180 0 0 VSS
port 1 nsew
flabel metal3 s 24732 70 24732 70 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 26970 70 26970 70 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 29213 70 29213 70 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 844 70 844 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 6958 70 6958 70 0 FreeSans 280 180 0 0 VSS
port 1 nsew
flabel metal3 s 14518 70 14518 70 0 FreeSans 280 180 0 0 VSS
port 1 nsew
flabel metal3 s 20167 70 20167 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 15687 70 15687 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 16527 70 16527 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 17437 70 17437 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 18347 70 18347 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 19257 70 19257 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 1777 70 1777 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 25571 70 25571 70 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 27809 70 27809 70 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 30053 70 30053 70 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 4439 70 4439 70 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 5279 70 5279 70 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 6119 70 6119 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 7799 70 7799 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 9060 70 9060 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 10319 70 10319 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 11999 70 11999 70 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 12839 70 12839 70 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 13679 70 13679 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 3600 70 3600 70 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 11160 70 11160 70 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 36213 70 36213 70 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 41200 70 41200 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 39380 70 39380 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 40290 70 40290 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 30893 70 30893 70 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 42110 70 42110 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 32573 70 32573 70 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 31733 70 31733 70 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 33413 70 33413 70 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 38470 70 38470 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 34346 70 34346 70 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 37085 70 37085 70 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 35263 70 35263 70 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal2 s 37718 70 37718 70 0 FreeSans 280 0 0 0 A[6]
port 4 nsew
flabel metal2 s 19633 70 19633 70 0 FreeSans 280 0 0 0 CLK
port 5 nsew
flabel metal2 s 1383 70 1383 70 0 FreeSans 280 0 0 0 D[0]
port 6 nsew
flabel metal2 s 21679 70 21679 70 0 FreeSans 280 0 0 0 A[2]
port 8 nsew
flabel metal2 s 22864 70 22864 70 0 FreeSans 280 0 0 0 A[1]
port 9 nsew
flabel metal2 s 24048 70 24048 70 0 FreeSans 280 0 0 0 A[0]
port 10 nsew
flabel metal2 s 9967 70 9967 70 0 FreeSans 280 180 0 0 Q[2]
port 11 nsew
flabel metal2 s 15673 70 15673 70 0 FreeSans 280 180 0 0 Q[3]
port 12 nsew
flabel metal2 s 35317 70 35317 70 0 FreeSans 280 0 0 0 CEN
port 13 nsew
flabel metal2 s 38170 70 38170 70 0 FreeSans 280 0 0 0 A[5]
port 14 nsew
flabel metal2 s 38693 70 38693 70 0 FreeSans 280 0 0 0 A[4]
port 15 nsew
flabel metal2 s 16461 70 16461 70 0 FreeSans 280 180 0 0 WEN[3]
port 16 nsew
flabel metal2 s 16734 70 16734 70 0 FreeSans 280 180 0 0 D[3]
port 19 nsew
flabel metal2 s 8622 70 8622 70 0 FreeSans 280 180 0 0 D[1]
port 20 nsew
flabel metal2 s 9496 70 9496 70 0 FreeSans 280 180 0 0 D[2]
port 21 nsew
flabel metal2 s 39463 70 39463 70 0 FreeSans 280 0 0 0 A[3]
port 22 nsew
flabel metal2 s 8151 70 8151 70 0 FreeSans 280 180 0 0 Q[1]
port 23 nsew
flabel metal2 s 9216 70 9216 70 0 FreeSans 280 180 0 0 WEN[2]
port 28 nsew
flabel metal2 s 8901 70 8901 70 0 FreeSans 280 180 0 0 WEN[1]
port 29 nsew
flabel metal2 s 28490 70 28490 70 0 FreeSans 280 0 0 0 GWEN
port 37 nsew
flabel metal3 s 59416 70 59416 70 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 43756 70 43756 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 57843 70 57843 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 42820 70 42820 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 56862 70 56862 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal2 s 58238 70 58238 70 0 FreeSans 280 180 0 0 D[7]
port 17 nsew
flabel metal2 s 57176 70 57176 70 0 FreeSans 280 180 0 0 Q[7]
port 18 nsew
flabel metal2 s 51470 70 51470 70 0 FreeSans 280 180 0 0 Q[6]
port 24 nsew
flabel metal2 s 43949 70 43949 70 0 FreeSans 280 180 0 0 Q[4]
port 26 nsew
flabel metal2 s 43358 70 43358 70 0 FreeSans 280 180 0 0 WEN[4]
port 30 nsew
flabel metal2 s 57764 70 57764 70 0 FreeSans 280 180 0 0 WEN[7]
port 31 nsew
flabel metal2 s 50719 70 50719 70 0 FreeSans 280 180 0 0 WEN[6]
port 32 nsew
flabel metal2 s 42891 70 42891 70 0 FreeSans 280 180 0 0 D[4]
port 33 nsew
flabel metal2 s 50999 70 50999 70 0 FreeSans 280 180 0 0 D[6]
port 34 nsew
flabel metal2 s 49925 70 49925 70 0 FreeSans 280 180 0 0 D[5]
port 25 nsew
flabel metal2 s 50204 70 50204 70 0 FreeSans 280 180 0 0 WEN[5]
port 27 nsew
flabel metal2 s 49454 70 49454 70 0 FreeSans 280 180 0 0 Q[5]
port 35 nsew
flabel metal3 s 55822 70 55822 70 0 FreeSans 280 180 0 0 VSS
port 1 nsew
flabel metal3 s 53302 70 53302 70 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 47422 70 47422 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 49102 70 49102 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 50361 70 50361 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 51622 70 51622 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 46582 70 46582 70 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 45742 70 45742 70 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 54982 70 54982 70 0 FreeSans 280 180 0 0 VDD
port 2 nsew
flabel metal3 s 54142 70 54142 70 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 48262 70 48262 70 0 FreeSans 280 180 0 0 VSS
port 1 nsew
flabel metal3 s 44902 70 44902 70 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 52462 70 52462 70 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal2 s 2844 70 2844 70 0 FreeSans 280 0 0 0 Q[0]
port 36 nsew
flabel metal2 s 2095 70 2095 70 0 FreeSans 280 0 0 0 WEN[0]
port 38 nsew
flabel metal3 s 31898 44921 31898 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 32769 44921 32769 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 40632 44921 40632 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 33626 44921 33626 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 37148 44921 37148 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 38333 44921 38333 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 34580 44921 34580 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 25140 44921 25140 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 7025 44921 7025 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 10805 44921 10805 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 4103 44921 4103 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 11663 44921 11663 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 3245 44921 3245 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 7883 44921 7883 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 27359 44921 27359 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 21847 44921 21847 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 14807 44921 14807 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 18950 44921 18950 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 29211 44921 29211 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 18110 44921 18110 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 16440 44921 16440 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 17298 44921 17298 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 13948 44921 13948 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 13090 44921 13090 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 1360 44921 1360 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 2218 44921 2218 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 10038 44921 10038 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 9180 44921 9180 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 20013 44921 20013 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 20991 44921 20991 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 30201 44921 30201 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 31099 44921 31099 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 28417 44921 28417 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 6128 44921 6128 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 5270 44921 5270 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 23166 44921 23166 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 24316 44921 24316 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 26363 44921 26363 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 35825 44921 35825 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 39693 44921 39693 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 49386 44921 49386 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 53166 44921 53166 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 54173 44921 54173 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 48529 44921 48529 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 52309 44921 52309 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 44749 44921 44749 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 59416 44921 59416 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 45606 44921 45606 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 55031 44921 55031 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 58371 44921 58371 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 57513 44921 57513 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 47221 44921 47221 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 46363 44921 46363 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 43311 44921 43311 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 42453 44921 42453 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 51121 44921 51121 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 50263 44921 50263 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal3 s 41453 44921 41453 44921 0 FreeSans 280 0 0 0 VSS
port 1 nsew
flabel metal3 s 56210 44921 56210 44921 0 FreeSans 280 0 0 0 VDD
port 2 nsew
flabel metal2 s 20870 70 20870 70 0 FreeSans 280 0 0 0 A[7]
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 60260 44986
string path 63.580 0.000 63.580 1.000 
<< end >>
