magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal2 >>
rect -119 704 119 732
rect -119 -704 -93 704
rect 93 -704 119 704
rect -119 -732 119 -704
<< via2 >>
rect -93 -704 93 704
<< metal3 >>
rect -119 704 119 732
rect -119 -704 -93 704
rect 93 -704 119 704
rect -119 -732 119 -704
<< end >>
