magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< psubdiff >>
rect -56 1737 56 1771
rect -56 -1737 -23 1737
rect 23 -1737 56 1737
rect -56 -1771 56 -1737
<< psubdiffcont >>
rect -23 -1737 23 1737
<< metal1 >>
rect -49 1737 49 1765
rect -49 -1737 -23 1737
rect 23 -1737 49 1737
rect -49 -1765 49 -1737
<< end >>
