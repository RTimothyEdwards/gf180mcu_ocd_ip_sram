magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -1782 158 1782 165
rect -1782 -158 -1775 158
rect 1775 -158 1782 158
rect -1782 -165 1782 -158
<< via2 >>
rect -1775 -158 1775 158
<< metal3 >>
rect -1782 158 1782 165
rect -1782 -158 -1775 158
rect 1775 -158 1782 158
rect -1782 -165 1782 -158
<< end >>
