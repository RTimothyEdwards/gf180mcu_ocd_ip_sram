magic
tech gf180mcuD
magscale 1 10
timestamp 1765482800
<< error_s >>
rect 19225 104090 19230 104095
rect 19271 25190 19276 104090
rect 39909 25190 39915 104095
rect 19209 23786 19236 23842
rect 19225 23780 19230 23786
rect 19265 23448 19292 23786
<< psubdiff >>
rect 18967 25183 20040 104192
rect 39151 25183 40172 104502
rect 59602 2309 59871 104499
<< metal1 >>
rect 0 2187 700 104470
<< metal2 >>
rect 296 2187 996 104477
<< metal3 >>
rect 296 2722 997 2791
rect 296 1905 996 2722
use M1_PSUB4310591302043_3v1024x8m81  M1_PSUB4310591302043_3v1024x8m81_0
timestamp 1764525316
transform -1 0 59970 0 1 104185
box 171 -29 59921 289
use M1_PSUB4310591302043_3v1024x8m81  M1_PSUB4310591302043_3v1024x8m81_1
timestamp 1764525316
transform -1 0 59970 0 1 2339
box 171 -29 59921 289
use M1_PSUB4310591302044_3v1024x8m81  M1_PSUB4310591302044_3v1024x8m81_0
timestamp 1765482800
transform 1 0 59631 0 1 798
box -29 1830 240 103358
use M1_PSUB4310591302044_3v1024x8m81  M1_PSUB4310591302044_3v1024x8m81_1
timestamp 1765482800
transform 1 0 18997 0 1 798
box -29 1830 240 103358
use M1_PSUB4310591302044_3v1024x8m81  M1_PSUB4310591302044_3v1024x8m81_2
timestamp 1765482800
transform 1 0 39932 0 1 798
box -29 1830 240 103358
use M1_PSUB4310591302044_3v1024x8m81  M1_PSUB4310591302044_3v1024x8m81_3
timestamp 1765482800
transform 1 0 78 0 1 798
box -29 1830 240 103358
use M1_PSUB4310591302045_3v1024x8m81  M1_PSUB4310591302045_3v1024x8m81_0
timestamp 1765482800
transform 1 0 39286 0 1 25213
box -29 -29 589 78883
use M1_PSUB4310591302045_3v1024x8m81  M1_PSUB4310591302045_3v1024x8m81_1
timestamp 1765482800
transform 1 0 19294 0 1 25213
box -29 -29 589 78883
use M1_PSUB4310591302046_3v1024x8m81  M1_PSUB4310591302046_3v1024x8m81_0
timestamp 1764525316
transform 1 0 19294 0 1 23477
box -29 -29 20539 309
<< labels >>
flabel metal3 s 646 2029 646 2029 0 FreeSans 313 0 0 0 VDD
port 1 nsew
<< properties >>
string path 4.620 11.160 4.620 0.000 
<< end >>
