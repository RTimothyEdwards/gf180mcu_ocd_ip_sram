magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< error_s >>
rect 9 -6018 48 -5962
rect 65 -6036 104 -6018
rect 138 -6036 177 -5962
<< nwell >>
rect -29 -1908 695 -1834
rect -30 -2230 695 -1908
<< nmos >>
rect 145 -5592 201 -4427
rect 305 -5592 361 -4427
rect 465 -5592 521 -4427
<< ndiff >>
rect 54 -4440 145 -4427
rect 54 -5567 70 -4440
rect 116 -5567 145 -4440
rect 54 -5592 145 -5567
rect 201 -5592 305 -4427
rect 361 -5592 465 -4427
rect 521 -4440 618 -4427
rect 521 -5567 550 -4440
rect 597 -5567 618 -4440
rect 521 -5592 618 -5567
<< ndiffc >>
rect 70 -5567 116 -4440
rect 550 -5567 597 -4440
<< psubdiff >>
rect 0 137 674 171
rect 0 91 141 137
rect 519 91 674 137
rect 0 56 674 91
rect 0 -5778 674 -5744
rect 0 -5824 141 -5778
rect 519 -5824 674 -5778
rect 0 -5859 674 -5824
<< nsubdiff >>
rect 0 -2057 670 -2025
rect 0 -2103 133 -2057
rect 401 -2103 670 -2057
rect 0 -2137 670 -2103
<< psubdiffcont >>
rect 141 91 519 137
rect 141 -5824 519 -5778
<< nsubdiffcont >>
rect 133 -2103 401 -2057
<< polysilicon >>
rect 145 -590 201 -558
rect 305 -590 361 -558
rect 465 -590 521 -558
rect 145 -686 521 -590
rect 145 -694 201 -686
rect 305 -694 361 -686
rect 465 -694 521 -686
rect 145 -1868 201 -1834
rect 305 -1868 361 -1834
rect 465 -1868 521 -1834
rect 137 -1963 535 -1868
rect 145 -4427 201 -3328
rect 305 -4427 361 -3328
rect 465 -4427 521 -3328
rect 145 -5643 201 -5592
rect 305 -5643 361 -5592
rect 465 -5643 521 -5592
<< metal1 >>
rect 0 137 674 165
rect 0 91 141 137
rect 519 91 674 137
rect 0 -38 674 91
rect 60 -39 142 -38
rect 60 -175 141 -39
rect 374 -175 455 -38
rect 217 -594 298 -465
rect 531 -594 611 -462
rect 217 -677 611 -594
rect 217 -778 298 -677
rect 531 -778 611 -677
rect 139 -1957 611 -1874
rect 0 -2057 455 -2039
rect 0 -2103 133 -2057
rect 401 -2103 455 -2057
rect 0 -2122 455 -2103
rect 55 -2191 137 -2122
rect 374 -2184 455 -2122
rect 531 -2366 611 -1957
rect -40 -3441 714 -3376
rect -40 -3582 714 -3518
rect -40 -3723 714 -3659
rect -40 -3864 714 -3800
rect -40 -4005 714 -3941
rect -40 -4147 714 -4082
rect 60 -4440 142 -4430
rect 60 -5567 70 -4440
rect 116 -5567 142 -4440
rect 60 -5648 142 -5567
rect 531 -4440 612 -4430
rect 531 -5567 550 -4440
rect 597 -5012 612 -4440
rect 597 -5567 611 -5012
rect 531 -5586 611 -5567
rect 56 -5649 146 -5648
rect 5 -5778 674 -5649
rect 5 -5824 141 -5778
rect 519 -5824 674 -5778
rect 5 -5852 674 -5824
<< metal2 >>
rect 147 -499 301 228
rect 49 -2178 137 -1710
rect 368 -2179 456 -1711
rect 213 -3284 616 -3038
rect 527 -4676 616 -3284
<< metal3 >>
rect -36 -647 774 -66
rect -40 -3464 774 -1981
rect 0 -5063 674 -4586
rect -46 -5510 774 -5144
use M1_POLY24310591302060_256x8m81  M1_POLY24310591302060_256x8m81_0
timestamp 1763766357
transform 1 0 343 0 1 -1914
box -128 -36 128 36
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_0
timestamp 1763766357
transform 1 0 571 0 1 -3161
box -43 -122 43 122
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_1
timestamp 1763766357
transform 1 0 258 0 1 -3161
box -43 -122 43 122
use M2_M1$$43376684_256x8m81  M2_M1$$43376684_256x8m81_0
timestamp 1763766357
transform 1 0 571 0 1 -5051
box -44 21 44 579
use M2_M1$$43379756_256x8m81  M2_M1$$43379756_256x8m81_0
timestamp 1763766357
transform 1 0 420 0 1 -230
box -44 -275 44 275
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_0
timestamp 1763766357
transform 1 0 93 0 1 -1528
box -44 -198 44 198
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_1
timestamp 1763766357
transform 1 0 415 0 1 -1528
box -44 -198 44 198
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_2
timestamp 1763766357
transform 1 0 256 0 1 -299
box -44 -198 44 198
use M2_M1$$47327276_256x8m81  M2_M1$$47327276_256x8m81_0
timestamp 1763766357
transform 1 0 93 0 1 -5505
box -45 -331 45 961
use M2_M1$$47515692_256x8m81  M2_M1$$47515692_256x8m81_0
timestamp 1763766357
transform 1 0 93 0 1 -2456
box -44 -504 44 284
use M2_M1$$47515692_256x8m81  M2_M1$$47515692_256x8m81_1
timestamp 1763766357
transform 1 0 93 0 1 -2456
box -44 -504 44 284
use M2_M1$$47515692_256x8m81  M2_M1$$47515692_256x8m81_2
timestamp 1763766357
transform 1 0 412 0 1 -2456
box -44 -504 44 284
use M2_M1$$47515692_256x8m81  M2_M1$$47515692_256x8m81_3
timestamp 1763766357
transform 1 0 412 0 1 -2456
box -44 -504 44 284
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_2
timestamp 1763766357
transform 1 0 93 0 1 -4743
box -45 -198 45 198
use M3_M2$$47332396_256x8m81  M3_M2$$47332396_256x8m81_0
timestamp 1763766357
transform 1 0 93 0 1 -2456
box -45 -504 45 504
use M3_M2$$47332396_256x8m81  M3_M2$$47332396_256x8m81_1
timestamp 1763766357
transform 1 0 93 0 1 -2456
box -45 -504 45 504
use M3_M2$$47332396_256x8m81  M3_M2$$47332396_256x8m81_2
timestamp 1763766357
transform 1 0 412 0 1 -2456
box -45 -504 45 504
use M3_M2$$47332396_256x8m81  M3_M2$$47332396_256x8m81_3
timestamp 1763766357
transform 1 0 412 0 1 -2456
box -45 -504 45 504
use M3_M2$$47333420_256x8m81  M3_M2$$47333420_256x8m81_0
timestamp 1763766357
transform 1 0 93 0 1 -5851
box -84 -185 84 275
use M3_M2$$47333420_256x8m81  M3_M2$$47333420_256x8m81_1
timestamp 1763766357
transform 1 0 420 0 1 -340
box -84 -185 84 275
use nmos_1p2$$47514668_256x8m81  nmos_1p2$$47514668_256x8m81_0
timestamp 1763766357
transform 1 0 159 0 -1 -95
box -102 -44 130 467
use nmos_1p2$$47514668_256x8m81  nmos_1p2$$47514668_256x8m81_1
timestamp 1763766357
transform 1 0 319 0 -1 -95
box -102 -44 130 467
use nmos_1p2$$47514668_256x8m81  nmos_1p2$$47514668_256x8m81_2
timestamp 1763766357
transform 1 0 479 0 -1 -95
box -102 -44 130 467
use pmos_1p2$$47512620_256x8m81  pmos_1p2$$47512620_256x8m81_0
timestamp 1763766357
transform 1 0 159 0 1 -3289
box -188 -86 216 1059
use pmos_1p2$$47512620_256x8m81  pmos_1p2$$47512620_256x8m81_1
timestamp 1763766357
transform 1 0 479 0 1 -3289
box -188 -86 216 1059
use pmos_1p2$$47512620_256x8m81  pmos_1p2$$47512620_256x8m81_3
timestamp 1763766357
transform 1 0 319 0 1 -3289
box -188 -86 216 1059
use pmos_1p2$$47513644_256x8m81  pmos_1p2$$47513644_256x8m81_0
timestamp 1763766357
transform 1 0 319 0 -1 -736
box -188 -86 216 1144
use pmos_1p2$$47513644_256x8m81  pmos_1p2$$47513644_256x8m81_1
timestamp 1763766357
transform 1 0 479 0 -1 -736
box -188 -86 216 1144
use pmos_1p2$$47513644_256x8m81  pmos_1p2$$47513644_256x8m81_2
timestamp 1763766357
transform 1 0 159 0 -1 -736
box -188 -86 216 1144
<< end >>
