magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< nmos >>
rect 0 0 56 246
<< ndiff >>
rect -88 233 0 246
rect -88 13 -75 233
rect -29 13 0 233
rect -88 0 0 13
rect 56 233 144 246
rect 56 13 85 233
rect 131 13 144 233
rect 56 0 144 13
<< ndiffc >>
rect -75 13 -29 233
rect 85 13 131 233
<< polysilicon >>
rect 0 246 56 291
rect 0 -44 56 0
<< metal1 >>
rect -75 233 -29 246
rect -75 0 -29 13
rect 85 233 131 246
rect 85 0 131 13
<< labels >>
flabel ndiffc -40 123 -40 123 0 FreeSans 93 0 0 0 S
flabel ndiffc 96 123 96 123 0 FreeSans 93 0 0 0 D
<< end >>
