magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal1 >>
rect -70 322 70 330
rect -70 -322 -61 322
rect 61 -322 70 322
rect -70 -330 70 -322
<< via1 >>
rect -61 -322 61 322
<< metal2 >>
rect -70 322 70 330
rect -70 -322 -61 322
rect 61 -322 70 322
rect -70 -330 70 -322
<< end >>
