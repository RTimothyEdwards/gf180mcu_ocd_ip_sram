magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -35 92 35 99
rect -35 -92 -28 92
rect 28 -92 35 92
rect -35 -99 35 -92
<< via2 >>
rect -28 -92 28 92
<< metal3 >>
rect -35 92 35 99
rect -35 -92 -28 92
rect 28 -92 35 92
rect -35 -99 35 -92
<< end >>
