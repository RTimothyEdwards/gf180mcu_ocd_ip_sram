magic
tech gf180mcuD
magscale 1 10
timestamp 1763585189
<< nwell >>
rect -371 3355 531 3507
rect -371 2774 3558 3355
rect -371 2024 3622 2774
rect -371 756 -57 819
rect 2474 756 2915 757
rect 3393 756 3622 795
rect -371 298 3622 756
rect -371 244 -44 298
<< polysilicon >>
rect 1589 3864 2442 3906
rect 116 3288 172 3616
rect 276 3288 332 3616
rect 753 3453 809 3475
rect 913 3453 969 3475
rect 1075 3453 1131 3475
rect 1235 3453 1291 3475
rect 1397 3453 1453 3460
rect 462 3411 1453 3453
rect 753 3190 809 3411
rect 913 3190 969 3411
rect 1074 3190 1130 3411
rect 1589 3340 1629 3864
rect 1742 3753 1798 3864
rect 1902 3753 1958 3864
rect 2064 3753 2120 3864
rect 2224 3753 2280 3864
rect 2386 3753 2442 3864
rect 2735 3383 2791 3468
rect 1234 3298 1629 3340
rect 1234 3190 1290 3298
rect 1409 3278 1629 3298
rect 1783 3331 2791 3383
rect 2895 3331 2951 3468
rect 3055 3331 3111 3468
rect 3215 3331 3271 3468
rect 1783 3288 3283 3331
rect 1409 3095 1572 3278
rect 1783 3155 1839 3288
rect 1943 3155 1999 3288
rect 2104 3155 2160 3288
rect 2264 3155 2320 3288
rect 2425 3155 2481 3288
rect 2585 3155 2641 3288
rect 2746 3155 2802 3288
rect 2906 3155 2962 3288
rect 3067 3155 3123 3288
rect 3227 3155 3283 3288
rect 116 2882 172 2893
rect 276 2882 332 2893
rect 116 2786 332 2882
rect 89 2094 145 2126
rect 249 2094 305 2126
rect 410 2094 466 2126
rect 570 2094 626 2126
rect 731 2094 787 2126
rect 891 2094 947 2126
rect 1052 2094 1108 2126
rect 1212 2094 1268 2126
rect 1373 2094 1429 2126
rect 1533 2094 1589 2126
rect 89 2051 1611 2094
rect 266 1850 322 2051
rect 428 1850 484 2051
rect 588 1850 644 2051
rect 750 1850 806 2051
rect 910 1850 966 2051
rect 1072 1850 1128 2051
rect 1232 2007 1611 2051
rect 1232 1850 1288 2007
rect 2010 1896 2066 2095
rect 1850 1850 2066 1896
rect 1906 1848 2066 1850
rect 2171 1848 2227 2095
rect 2331 1848 2387 2095
rect 2636 2065 2692 2097
rect 2501 2063 2692 2065
rect 2797 2063 2853 2097
rect 2501 2060 2856 2063
rect 2957 2060 3013 2095
rect 2501 2017 3013 2060
rect 2501 2007 2856 2017
rect 1906 1840 2010 1848
rect 2640 1847 2696 2007
rect 2800 1847 2856 2007
rect 1689 1423 1745 1550
rect 2171 1423 2227 1549
rect 1689 1381 2227 1423
rect 122 1200 810 1201
rect 115 1199 810 1200
rect 115 1158 813 1199
rect 115 1067 171 1158
rect 275 1067 331 1158
rect 436 1067 492 1158
rect 596 1067 652 1158
rect 757 1067 813 1158
rect 115 850 171 899
rect 275 850 331 899
rect 436 850 492 899
rect 596 850 652 899
rect 757 850 813 899
rect 115 753 186 850
rect 275 753 346 850
rect 436 753 507 850
rect 596 753 667 850
rect 757 753 828 850
rect 1149 849 1209 904
rect 940 790 1209 849
rect 130 656 186 753
rect 290 656 346 753
rect 451 656 507 753
rect 611 656 667 753
rect 772 656 828 753
rect 1153 675 1209 790
rect 1313 675 1369 898
rect 1656 890 1716 897
rect 1447 831 1716 890
rect 1660 679 1716 831
rect 1820 679 1876 897
rect 2153 847 2209 899
rect 1957 789 2213 847
rect 2321 815 2377 899
rect 2653 847 2709 898
rect 2157 678 2213 789
rect 2317 678 2373 815
rect 2446 789 2709 847
rect 2985 819 3041 853
rect 2653 703 2709 789
rect 2931 760 2975 819
rect 2985 760 3202 819
rect 2985 658 3041 760
rect 3145 656 3201 760
<< metal1 >>
rect 833 3871 2517 3917
rect 833 3815 913 3871
rect 201 3584 248 3749
rect 832 3687 913 3815
rect 1144 3601 1225 3871
rect 1458 3601 1539 3871
rect 1827 3601 1873 3871
rect 2149 3597 2195 3871
rect 2471 3659 2517 3871
rect 2804 3857 3198 3906
rect 201 3531 534 3584
rect 201 3236 248 3531
rect 483 3363 534 3531
rect 1667 3390 1713 3574
rect 1988 3390 2034 3572
rect 2310 3390 2356 3587
rect 830 3306 2356 3390
rect 830 3136 912 3306
rect 1144 3127 1225 3306
rect 2288 3294 2356 3306
rect 2288 3293 2345 3294
rect 1865 2812 1946 3050
rect 2177 2812 2258 3065
rect 2491 2812 2572 3065
rect 2804 2812 2886 3857
rect 3117 2812 3198 3857
rect 184 2747 729 2800
rect 1865 2744 3198 2812
rect 37 2604 1688 2688
rect 37 2327 119 2604
rect 323 2355 404 2604
rect 637 2355 717 2604
rect 981 2355 1062 2604
rect 1283 2355 1364 2604
rect 1607 2430 1688 2604
rect 166 2083 247 2251
rect 490 2083 570 2232
rect 813 2083 894 2220
rect 1136 2083 1218 2213
rect 166 2073 1218 2083
rect 1450 2073 1531 2335
rect 166 1999 1531 2073
rect 1605 2008 1814 2093
rect 2077 2086 2158 2211
rect 2415 2086 2474 2196
rect 1920 2003 2558 2086
rect 166 1740 247 1999
rect 490 1740 570 1999
rect 813 1740 894 1999
rect 1136 1740 1218 1999
rect 353 1553 434 1740
rect 667 1553 747 1740
rect 980 1553 1061 1740
rect 1309 1553 1359 1634
rect 1920 1556 2002 2003
rect 2704 1723 2786 2206
rect 3024 2002 3100 2217
rect 353 1501 1359 1553
rect 604 1377 3129 1445
rect 3201 1293 3468 1518
rect -261 1197 3517 1293
rect 851 1060 1122 1128
rect 211 853 260 1000
rect 536 853 585 1000
rect 851 853 900 1060
rect 1070 897 1124 987
rect 1293 941 1341 1132
rect 211 770 989 853
rect 211 551 260 770
rect 512 769 585 770
rect 826 769 900 770
rect 536 543 585 769
rect 854 553 900 769
rect 1078 568 1124 897
rect 1287 891 1347 941
rect 1400 938 1476 1022
rect 1293 841 1341 891
rect 1425 568 1476 938
rect 1559 842 1610 1004
rect 1559 794 1848 842
rect 1559 568 1610 794
rect 1933 568 1983 1004
rect 2065 842 2116 1004
rect 2406 920 2499 1004
rect 2065 794 2355 842
rect 2065 562 2116 794
rect 2452 695 2499 920
rect 2421 562 2499 695
rect 2578 554 2625 993
rect 2593 553 2625 554
rect 3070 457 3120 1005
<< metal2 >>
rect 602 1377 667 2816
rect 1437 2663 1502 3231
rect 1592 2797 1654 3383
rect 1592 2733 2006 2797
rect 1437 2595 1879 2663
rect 1943 2604 2006 2733
rect 1813 1950 1879 2595
rect 1144 1882 2296 1950
rect 1144 1066 1210 1882
rect 3063 863 3129 1445
rect 3201 1199 3468 1518
rect 1052 754 2792 821
<< metal3 >>
rect -250 3588 3587 3958
rect -252 2173 3500 3126
rect 2712 2088 2779 2089
rect 3028 2088 3093 2089
rect 1532 2021 3093 2088
rect -252 1592 3500 1952
rect -261 1187 3517 1528
rect -252 822 3500 1125
rect -252 408 3514 726
use M1_NWELL02_512x8m81  M1_NWELL02_512x8m81_0
timestamp 1763564386
transform 1 0 -217 0 -1 575
box -154 -159 154 159
use M1_NWELL03_512x8m81  M1_NWELL03_512x8m81_0
timestamp 1763564386
transform 1 0 3413 0 1 2329
box -210 -445 210 445
use M1_NWELL04_512x8m81  M1_NWELL04_512x8m81_0
timestamp 1763564386
transform 1 0 -217 0 1 2329
box -154 -445 154 445
use M1_PACTIVE4310591302034_512x8m81  M1_PACTIVE4310591302034_512x8m81_0
timestamp 1763564386
transform 1 0 -217 0 1 3762
box -36 -128 36 128
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_0
timestamp 1763564386
transform 1 0 688 0 1 1239
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_1
timestamp 1763564386
transform 1 0 240 0 1 1239
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_2
timestamp 1763564386
transform 1 0 224 0 1 2834
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_3
timestamp 1763564386
transform 1 0 530 0 1 3405
box -67 -48 67 47
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_0
timestamp 1763564386
transform -1 0 1476 0 1 3151
box -96 -124 67 124
use M1_POLY2$$45109292_512x8m81  M1_POLY2$$45109292_512x8m81_0
timestamp 1763564386
transform 1 0 2073 0 1 3335
box -289 -48 289 48
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1763564386
transform 1 0 2475 0 1 818
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1763564386
transform 1 0 2961 0 1 789
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_2
timestamp 1763564386
transform 1 0 2348 0 1 1908
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_3
timestamp 1763564386
transform 1 0 2527 0 1 2036
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_4
timestamp 1763564386
transform 1 0 1824 0 1 818
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_5
timestamp 1763564386
transform 1 0 1986 0 1 818
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_6
timestamp 1763564386
transform 1 0 2331 0 1 818
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_7
timestamp 1763564386
transform 1 0 1459 0 1 861
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_8
timestamp 1763564386
transform 1 0 942 0 1 819
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_9
timestamp 1763564386
transform 1 0 1560 0 1 1895
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_10
timestamp 1763564386
transform 1 0 1317 0 1 861
box -36 -36 36 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_0
timestamp 1763564386
transform 1 0 2019 0 1 2635
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_1
timestamp 1763564386
transform 1 0 1671 0 1 2056
box -62 -36 62 36
use M1_PSUB$$44997676_512x8m81  M1_PSUB$$44997676_512x8m81_0
timestamp 1763564386
transform 1 0 3357 0 -1 1700
box -165 -114 166 114
use M1_PSUB$$44997676_512x8m81  M1_PSUB$$44997676_512x8m81_1
timestamp 1763564386
transform 1 0 -106 0 -1 1700
box -165 -114 166 114
use M1_PSUB_285_512x8m81  M1_PSUB_285_512x8m81_0
timestamp 1763564386
transform 1 0 3413 0 -1 1065
box -118 -58 111 57
use M1_PSUB_285_512x8m81  M1_PSUB_285_512x8m81_1
timestamp 1763564386
transform 1 0 -171 0 -1 1065
box -118 -58 111 57
use M2_M1$$43374636_512x8m81  M2_M1$$43374636_512x8m81_0
timestamp 1763564386
transform 1 0 170 0 1 1323
box -119 -123 119 123
use M2_M1$$45002796_512x8m81  M2_M1$$45002796_512x8m81_0
timestamp 1763564386
transform 1 0 2144 0 1 1246
box -783 -46 783 46
use M2_M1$$45003820_512x8m81  M2_M1$$45003820_512x8m81_0
timestamp 1763564386
transform 1 0 3320 0 1 1399
box -119 -198 119 128
use M2_M1c$$203396140_512x8m81  M2_M1c$$203396140_512x8m81_0
timestamp 1763564386
transform 1 0 697 0 1 2781
box -108 -46 108 46
use M3_M2$$45005868_512x8m81  M3_M2$$45005868_512x8m81_0
timestamp 1763564386
transform 1 0 2144 0 1 1246
box -783 -46 783 46
use M3_M2$$45006892_512x8m81  M3_M2$$45006892_512x8m81_0
timestamp 1763564386
transform 1 0 3320 0 1 1399
box -119 -198 119 118
use M3_M2$$45008940_512x8m81  M3_M2$$45008940_512x8m81_0
timestamp 1763564386
transform 1 0 170 0 1 1323
box -119 -123 119 123
use nmos_1p2$$45100076_512x8m81  nmos_1p2$$45100076_512x8m81_0
timestamp 1763564386
transform -1 0 2814 0 -1 1820
box -130 -44 263 287
use nmos_1p2$$45101100_512x8m81  nmos_1p2$$45101100_512x8m81_0
timestamp 1763564386
transform 1 0 241 0 1 918
box -214 -44 660 150
use nmos_1p2$$45102124_512x8m81  nmos_1p2$$45102124_512x8m81_0
timestamp 1763564386
transform -1 0 1106 0 -1 1820
box -270 -44 928 255
use nmos_1p2$$45103148_512x8m81  nmos_1p2$$45103148_512x8m81_0
timestamp 1763564386
transform -1 0 2233 0 -1 1820
box -242 -44 792 310
use nmos_5p04310591302012_512x8m81  nmos_5p04310591302012_512x8m81_0
timestamp 1763564386
transform -1 0 3188 0 1 3504
box -171 -44 541 255
use nmos_5p04310591302023_512x8m81  nmos_5p04310591302023_512x8m81_0
timestamp 1763564386
transform 1 0 2185 0 1 938
box -124 -44 285 100
use nmos_5p04310591302023_512x8m81  nmos_5p04310591302023_512x8m81_1
timestamp 1763564386
transform 1 0 1181 0 1 938
box -124 -44 285 100
use nmos_5p04310591302023_512x8m81  nmos_5p04310591302023_512x8m81_2
timestamp 1763564386
transform 1 0 1688 0 1 938
box -124 -44 285 100
use nmos_5p04310591302028_512x8m81  nmos_5p04310591302028_512x8m81_0
timestamp 1763564386
transform 1 0 849 0 1 3504
box -184 -44 692 255
use nmos_5p04310591302028_512x8m81  nmos_5p04310591302028_512x8m81_1
timestamp 1763564386
transform 1 0 1838 0 1 3504
box -184 -44 692 255
use nmos_5p04310591302032_512x8m81  nmos_5p04310591302032_512x8m81_0
timestamp 1763564386
transform -1 0 304 0 1 3656
box -116 -44 277 150
use nmos_5p04310591302033_512x8m81  nmos_5p04310591302033_512x8m81_0
timestamp 1763564386
transform 1 0 2653 0 1 938
box -92 -44 148 100
use nmos_5p04310591302034_512x8m81  nmos_5p04310591302034_512x8m81_0
timestamp 1763564386
transform 1 0 2985 0 1 892
box -88 -44 144 178
use pmos_1p2$$45095980_512x8m81  pmos_1p2$$45095980_512x8m81_0
timestamp 1763564386
transform -1 0 3017 0 1 2863
box -440 -86 1408 339
use pmos_1p2$$46281772_512x8m81  pmos_1p2$$46281772_512x8m81_0
timestamp 1763564386
transform -1 0 2943 0 -1 2555
box -244 -86 481 509
use pmos_1p2$$46281772_512x8m81  pmos_1p2$$46281772_512x8m81_1
timestamp 1763564386
transform -1 0 2317 0 -1 2555
box -244 -86 481 509
use pmos_1p2$$46282796_512x8m81  pmos_1p2$$46282796_512x8m81_0
timestamp 1763564386
transform 1 0 256 0 1 402
box -300 -86 746 297
use pmos_1p2$$46283820_512x8m81  pmos_1p2$$46283820_512x8m81_0
timestamp 1763564386
transform -1 0 1323 0 -1 2540
box -440 -86 1408 467
use pmos_1p2$$46284844_512x8m81  pmos_1p2$$46284844_512x8m81_0
timestamp 1763564386
transform 1 0 3027 0 1 457
box -216 -86 348 245
use pmos_1p2$$46285868_512x8m81  pmos_1p2$$46285868_512x8m81_0
timestamp 1763564386
transform 1 0 1248 0 1 2938
box -188 -86 216 297
use pmos_1p2$$46286892_512x8m81  pmos_1p2$$46286892_512x8m81_0
timestamp 1763564386
transform 1 0 823 0 1 2938
box -244 -86 481 297
use pmos_1p2$$46287916_512x8m81  pmos_1p2$$46287916_512x8m81_0
timestamp 1763564386
transform -1 0 290 0 1 2932
box -216 -86 348 404
use pmos_5p04310591302027_512x8m81  pmos_5p04310591302027_512x8m81_0
timestamp 1763564386
transform 1 0 2185 0 1 527
box -202 -86 362 198
use pmos_5p04310591302027_512x8m81  pmos_5p04310591302027_512x8m81_1
timestamp 1763564386
transform 1 0 1181 0 1 527
box -202 -86 362 198
use pmos_5p04310591302027_512x8m81  pmos_5p04310591302027_512x8m81_2
timestamp 1763564386
transform 1 0 1688 0 1 527
box -202 -86 362 198
use pmos_5p04310591302038_512x8m81  pmos_5p04310591302038_512x8m81_0
timestamp 1763564386
transform 1 0 2653 0 1 553
box -174 -86 230 198
use po_m1_512x8m81  po_m1_512x8m81_0
timestamp 1763564386
transform 1 0 1920 0 1 1328
box -21 0 113 95
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_0
timestamp 1763564386
transform 1 0 2232 0 1 408
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_1
timestamp 1763564386
transform 1 0 1726 0 1 408
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_2
timestamp 1763564386
transform -1 0 2465 0 -1 1805
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_3
timestamp 1763564386
transform 1 0 3436 0 1 901
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_4
timestamp 1763564386
transform 1 0 3436 0 1 1593
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_5
timestamp 1763564386
transform 1 0 3220 0 1 408
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_6
timestamp 1763564386
transform 1 0 2903 0 1 408
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_7
timestamp 1763564386
transform 1 0 2759 0 1 408
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_8
timestamp 1763564386
transform -1 0 2933 0 -1 1805
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_9
timestamp 1763564386
transform -1 0 2620 0 -1 1805
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_10
timestamp 1763564386
transform -1 0 1521 0 -1 1805
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_11
timestamp 1763564386
transform 1 0 50 0 1 455
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_12
timestamp 1763564386
transform -1 0 -184 0 -1 708
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_13
timestamp 1763564386
transform -1 0 1052 0 -1 1807
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_14
timestamp 1763564386
transform 1 0 -249 0 1 901
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_15
timestamp 1763564386
transform 1 0 -249 0 1 1593
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_16
timestamp 1763564386
transform 1 0 1218 0 1 408
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_17
timestamp 1763564386
transform 1 0 677 0 1 453
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_18
timestamp 1763564386
transform 1 0 364 0 1 454
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_19
timestamp 1763564386
transform 1 0 -249 0 1 2174
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_20
timestamp 1763564386
transform -1 0 79 0 -1 3871
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_21
timestamp 1763564386
transform -1 0 84 0 -1 3086
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_22
timestamp 1763564386
transform -1 0 745 0 -1 3811
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_23
timestamp 1763564386
transform -1 0 1052 0 -1 3811
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_24
timestamp 1763564386
transform -1 0 1379 0 -1 3811
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_25
timestamp 1763564386
transform -1 0 420 0 -1 3871
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_26
timestamp 1763564386
transform -1 0 408 0 -1 3086
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_27
timestamp 1763564386
transform -1 0 746 0 -1 3116
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_28
timestamp 1763564386
transform -1 0 1054 0 -1 3086
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_29
timestamp 1763564386
transform -1 0 83 0 -1 2545
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_30
timestamp 1763564386
transform -1 0 1054 0 -1 2545
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_31
timestamp 1763564386
transform -1 0 -184 0 -1 3885
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_32
timestamp 1763564386
transform -1 0 1359 0 -1 3086
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_33
timestamp 1763564386
transform 1 0 -249 0 1 2578
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_34
timestamp 1763564386
transform 1 0 3436 0 1 2174
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_35
timestamp 1763564386
transform 1 0 3436 0 1 2501
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_36
timestamp 1763564386
transform -1 0 2619 0 -1 2502
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_37
timestamp 1763564386
transform -1 0 2934 0 -1 2502
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_38
timestamp 1763564386
transform -1 0 2308 0 -1 2502
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_39
timestamp 1763564386
transform -1 0 2007 0 -1 2502
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_40
timestamp 1763564386
transform -1 0 1789 0 -1 3103
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_41
timestamp 1763564386
transform -1 0 2095 0 -1 3103
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_42
timestamp 1763564386
transform -1 0 2404 0 -1 3103
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_43
timestamp 1763564386
transform -1 0 2722 0 -1 3103
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_44
timestamp 1763564386
transform -1 0 3034 0 -1 3103
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_45
timestamp 1763564386
transform -1 0 3348 0 -1 3103
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_46
timestamp 1763564386
transform -1 0 2720 0 -1 3811
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_47
timestamp 1763564386
transform -1 0 3033 0 -1 3811
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_48
timestamp 1763564386
transform -1 0 3349 0 -1 3811
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_49
timestamp 1763564386
transform 0 -1 3198 1 0 2023
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_50
timestamp 1763564386
transform 0 -1 2848 1 0 2021
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_51
timestamp 1763564386
transform -1 0 1672 0 -1 2515
box -9 0 73 215
use via1_R90_512x8m81  via1_R90_512x8m81_0
timestamp 1763564386
transform 0 -1 1695 1 0 2022
box 0 0 65 89
use via1_x2_512x8m81  via1_x2_512x8m81_0
timestamp 1763564386
transform 1 0 1736 0 1 910
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_1
timestamp 1763564386
transform 1 0 2242 0 1 910
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_2
timestamp 1763564386
transform 1 0 2750 0 1 910
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_3
timestamp 1763564386
transform 1 0 2907 0 1 910
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_4
timestamp 1763564386
transform 1 0 3063 0 1 862
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_5
timestamp 1763564386
transform 1 0 1052 0 1 675
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_6
timestamp 1763564386
transform 1 0 1274 0 1 910
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_7
timestamp 1763564386
transform 1 0 50 0 1 910
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_8
timestamp 1763564386
transform 1 0 344 0 1 910
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_9
timestamp 1763564386
transform 1 0 674 0 1 910
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_10
timestamp 1763564386
transform -1 0 1501 0 -1 3231
box -8 0 72 222
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_0
timestamp 1763564386
transform 0 -1 3128 1 0 1378
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_1
timestamp 1763564386
transform 0 -1 3000 1 0 754
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_2
timestamp 1763564386
transform 0 -1 812 1 0 1378
box -8 0 72 215
use via1_x2_R270_512x8m81  via1_x2_R270_512x8m81_0
timestamp 1763564386
transform 0 1 2158 -1 0 1944
box -8 0 75 215
use via1_x2_R270_512x8m81  via1_x2_R270_512x8m81_1
timestamp 1763564386
transform 0 1 994 -1 0 1127
box -8 0 75 215
use via1_x2_R270_512x8m81  via1_x2_R270_512x8m81_2
timestamp 1763564386
transform 0 1 1944 -1 0 2676
box -8 0 75 215
use via1_x2_R270_512x8m81  via1_x2_R270_512x8m81_3
timestamp 1763564386
transform 0 1 1526 -1 0 1941
box -8 0 75 215
use via1_x2_R270_512x8m81  via1_x2_R270_512x8m81_4
timestamp 1763564386
transform 0 1 1592 -1 0 3383
box -8 0 75 215
use via2_x2_512x8m81  via2_x2_512x8m81_0
timestamp 1763564386
transform 1 0 2242 0 1 902
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_1
timestamp 1763564386
transform 1 0 1736 0 1 902
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_2
timestamp 1763564386
transform 1 0 2750 0 1 902
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_3
timestamp 1763564386
transform 1 0 2907 0 1 902
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_4
timestamp 1763564386
transform 1 0 674 0 1 902
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_5
timestamp 1763564386
transform 1 0 344 0 1 902
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_6
timestamp 1763564386
transform 1 0 50 0 1 902
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_7
timestamp 1763564386
transform 1 0 1274 0 1 902
box -9 0 74 222
use via2_x2_R90_512x8m81  via2_x2_R90_512x8m81_0
timestamp 1763564386
transform 0 -1 1747 1 0 2022
box -9 0 73 215
<< labels >>
rlabel metal3 s 1678 2661 1678 2661 4 vdd
port 1 nsew
rlabel metal3 s 1514 3810 1514 3810 4 vss
port 2 nsew
rlabel metal1 s 2846 3895 2846 3895 4 se
port 5 nsew
rlabel metal1 s 1019 2048 1019 2048 4 pcb
port 4 nsew
rlabel metal3 s 173 1495 173 1495 4 men
port 3 nsew
rlabel metal3 s 1601 1885 1601 1885 4 vss
port 2 nsew
rlabel metal3 s 1601 1812 1601 1812 4 vss
port 2 nsew
rlabel metal3 s 1042 705 1042 705 4 vdd
port 1 nsew
<< properties >>
string path 20.320 27.120 20.320 27.785 22.565 27.785 22.565 26.905 
<< end >>
