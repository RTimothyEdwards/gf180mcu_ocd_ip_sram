magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< polysilicon >>
rect -41 243 14 277
rect 118 243 173 277
rect -41 -34 14 0
rect 118 -34 173 0
use nmos_5p04310591302029_512x8m81  nmos_5p04310591302029_512x8m81_0
timestamp 1763476864
transform 1 0 -14 0 1 0
box -116 -44 277 287
<< end >>
