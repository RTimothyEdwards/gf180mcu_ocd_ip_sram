magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< error_p >>
rect -75 0 -29 84
rect 85 0 131 84
<< nwell >>
rect -174 -86 230 170
<< pmos >>
rect 0 0 56 84
<< pdiff >>
rect -88 71 0 84
rect -88 13 -75 71
rect -29 13 0 71
rect -88 0 0 13
rect 56 71 144 84
rect 56 13 85 71
rect 131 13 144 71
rect 56 0 144 13
<< pdiffc >>
rect -75 13 -29 71
rect 85 13 131 71
<< polysilicon >>
rect 0 84 56 128
rect 0 -44 56 0
<< metal1 >>
rect -75 71 -29 84
rect -75 0 -29 13
rect 85 71 131 84
rect 85 0 131 13
<< labels >>
flabel pdiffc -40 42 -40 42 0 FreeSans 186 0 0 0 S
flabel pdiffc 96 42 96 42 0 FreeSans 186 0 0 0 D
<< end >>
