magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< error_s >>
rect 911 2819 935 3075
<< nwell >>
rect 107 4947 1143 5223
rect 854 2649 935 4239
<< nmos >>
rect 483 911 539 2055
rect 612 911 668 2055
<< ndiff >>
rect 373 2031 483 2055
rect 373 1023 396 2031
rect 442 1023 483 2031
rect 373 911 483 1023
rect 539 911 612 2055
rect 668 2030 779 2055
rect 668 1023 710 2030
rect 756 1023 779 2030
rect 668 911 779 1023
<< ndiffc >>
rect 396 1023 442 2031
rect 710 1023 756 2030
<< psubdiff >>
rect 889 2020 982 2055
rect 889 375 911 2020
rect 959 375 982 2020
rect 889 340 982 375
rect 288 159 1009 184
rect 288 113 338 159
rect 847 113 1009 159
rect 288 88 1009 113
<< nsubdiff >>
rect 206 5074 1043 5107
rect 206 5028 320 5074
rect 436 5028 720 5074
rect 867 5028 1043 5074
rect 206 4995 1043 5028
<< psubdiffcont >>
rect 911 375 959 2020
rect 338 113 847 159
<< nsubdiffcont >>
rect 320 5028 436 5074
rect 720 5028 867 5074
<< polysilicon >>
rect 347 7027 403 7265
rect 507 7027 563 7265
rect 667 7027 723 7265
rect 827 7027 883 7265
rect 347 6954 883 7027
rect 347 6937 403 6954
rect 507 6937 563 6954
rect 667 6937 723 6954
rect 827 6937 883 6954
rect 347 5263 403 5801
rect 507 5263 563 5801
rect 667 5263 723 5801
rect 827 5263 883 5801
rect 345 5168 899 5263
rect 472 2656 528 2709
rect 472 2560 539 2656
rect 483 2055 539 2560
rect 632 2415 688 2709
rect 612 2347 688 2415
rect 612 2055 668 2347
rect 483 860 539 911
rect 612 860 668 911
<< metal1 >>
rect 268 7922 474 7982
rect 268 7646 349 7922
rect 581 7646 662 7980
rect 895 7646 976 7980
rect 416 7035 498 7366
rect 738 7035 819 7126
rect 416 6951 819 7035
rect 416 6846 498 6951
rect 738 6846 819 6951
rect 346 5174 898 5257
rect 535 5173 617 5174
rect 170 5074 459 5092
rect 170 5028 320 5074
rect 436 5028 459 5074
rect 170 5009 459 5028
rect 378 5008 459 5009
rect 378 4778 460 5008
rect 535 2730 616 5173
rect 692 5074 1043 5092
rect 692 5028 720 5074
rect 867 5028 1043 5074
rect 692 5009 1043 5028
rect 692 2741 976 5009
rect 255 2573 1068 2637
rect 255 2431 1068 2496
rect 255 2291 1068 2355
rect 255 2149 1068 2214
rect 378 2031 459 2048
rect 378 1023 396 2031
rect 442 1023 459 2031
rect 378 917 459 1023
rect 692 2030 976 2048
rect 692 1023 710 2030
rect 756 2020 976 2030
rect 756 1023 911 2020
rect 692 375 911 1023
rect 959 375 976 2020
rect 692 188 976 375
rect 692 181 981 188
rect 288 159 1009 181
rect 288 113 338 159
rect 847 113 1009 159
rect 288 91 1009 113
<< metal2 >>
rect 734 7097 889 7809
rect 692 3574 981 5058
rect 374 2741 620 2986
rect 374 1806 464 2741
rect 692 29 981 2048
<< metal3 >>
rect 107 7657 1038 7658
rect 107 6991 1039 7657
rect 107 6414 1038 6913
rect 107 5683 1036 6320
rect 107 3541 1036 5447
rect 598 1540 1038 2017
rect 598 730 1039 1366
rect 598 -24 1041 611
use M1_NACTIVE4310591302024_512x8m81  M1_NACTIVE4310591302024_512x8m81_0
timestamp 1763476864
transform 1 0 936 0 1 2947
box -38 -128 36 128
use M1_POLY24310591302059_512x8m81  M1_POLY24310591302059_512x8m81_0
timestamp 1763476864
transform 1 0 605 0 1 5215
box -161 -36 161 36
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1763476864
transform -1 0 576 0 1 2864
box -43 -122 43 122
use M2_M1$$43376684_512x8m81  M2_M1$$43376684_512x8m81_0
timestamp 1763476864
transform -1 0 419 0 1 1469
box -44 -579 44 579
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_0
timestamp 1763476864
transform 1 0 779 0 1 7372
box -44 -275 44 275
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_1
timestamp 1763476864
transform 1 0 616 0 1 7372
box -44 -275 44 275
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_2
timestamp 1763476864
transform -1 0 295 0 1 7372
box -44 -275 44 275
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_0
timestamp 1763476864
transform -1 0 295 0 1 6645
box -44 -198 44 198
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_1
timestamp 1763476864
transform 1 0 622 0 1 6645
box -44 -198 44 198
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_2
timestamp 1763476864
transform 1 0 935 0 1 6645
box -44 -198 44 198
use M2_M1$$47500332_512x8m81  M2_M1$$47500332_512x8m81_0
timestamp 1763476864
transform 1 0 737 0 1 4307
box -44 -732 44 732
use M2_M1$$47500332_512x8m81  M2_M1$$47500332_512x8m81_1
timestamp 1763476864
transform 1 0 421 0 1 4307
box -44 -732 44 732
use M2_M1$$47500332_512x8m81  M2_M1$$47500332_512x8m81_2
timestamp 1763476864
transform 1 0 935 0 1 4307
box -44 -732 44 732
use M2_M1$$47640620_512x8m81  M2_M1$$47640620_512x8m81_0
timestamp 1763476864
transform 1 0 935 0 1 1068
box -45 -884 45 884
use M2_M1$$47640620_512x8m81  M2_M1$$47640620_512x8m81_1
timestamp 1763476864
transform 1 0 737 0 1 1068
box -45 -884 45 884
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_0
timestamp 1763476864
transform 1 0 935 0 1 1753
box -45 -198 45 198
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_1
timestamp 1763476864
transform 1 0 737 0 1 1753
box -45 -198 45 198
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_2
timestamp 1763476864
transform -1 0 295 0 1 6645
box -45 -198 45 198
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_3
timestamp 1763476864
transform 1 0 622 0 1 6645
box -45 -198 45 198
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_4
timestamp 1763476864
transform 1 0 935 0 1 6645
box -45 -198 45 198
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_0
timestamp 1763476864
transform 1 0 935 0 1 306
box -45 -275 45 275
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_1
timestamp 1763476864
transform 1 0 737 0 1 306
box -45 -275 45 275
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_2
timestamp 1763476864
transform 1 0 616 0 1 7372
box -45 -275 45 275
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_3
timestamp 1763476864
transform -1 0 295 0 1 7372
box -45 -275 45 275
use M3_M2$$47644716_512x8m81  M3_M2$$47644716_512x8m81_0
timestamp 1763476864
transform 1 0 737 0 1 4307
box -45 -732 45 732
use M3_M2$$47644716_512x8m81  M3_M2$$47644716_512x8m81_1
timestamp 1763476864
transform 1 0 421 0 1 4307
box -45 -732 45 732
use M3_M2$$47644716_512x8m81  M3_M2$$47644716_512x8m81_2
timestamp 1763476864
transform 1 0 935 0 1 4307
box -45 -732 45 732
use nmos_1p2$$47641644_512x8m81  nmos_1p2$$47641644_512x8m81_0
timestamp 1763476864
transform -1 0 869 0 -1 7726
box -102 -44 130 467
use nmos_1p2$$47641644_512x8m81  nmos_1p2$$47641644_512x8m81_1
timestamp 1763476864
transform -1 0 549 0 -1 7726
box -102 -44 130 467
use nmos_1p2$$47641644_512x8m81  nmos_1p2$$47641644_512x8m81_2
timestamp 1763476864
transform -1 0 389 0 -1 7726
box -102 -44 130 467
use nmos_1p2$$47641644_512x8m81  nmos_1p2$$47641644_512x8m81_3
timestamp 1763476864
transform -1 0 709 0 -1 7726
box -102 -44 130 467
use pmos_1p2$$47513644_512x8m81  pmos_1p2$$47513644_512x8m81_0
timestamp 1763476864
transform -1 0 709 0 -1 6895
box -188 -86 216 1144
use pmos_1p2$$47513644_512x8m81  pmos_1p2$$47513644_512x8m81_1
timestamp 1763476864
transform -1 0 549 0 -1 6895
box -188 -86 216 1144
use pmos_1p2$$47513644_512x8m81  pmos_1p2$$47513644_512x8m81_2
timestamp 1763476864
transform -1 0 389 0 -1 6895
box -188 -86 216 1144
use pmos_1p2$$47513644_512x8m81  pmos_1p2$$47513644_512x8m81_3
timestamp 1763476864
transform -1 0 869 0 -1 6895
box -188 -86 216 1144
use pmos_1p2$$47642668_512x8m81  pmos_1p2$$47642668_512x8m81_0
timestamp 1763476864
transform -1 0 674 0 1 2735
box -194 -86 220 1504
use pmos_1p2$$47643692_512x8m81  pmos_1p2$$47643692_512x8m81_0
timestamp 1763476864
transform -1 0 514 0 1 2735
box -188 -86 216 1504
<< end >>
