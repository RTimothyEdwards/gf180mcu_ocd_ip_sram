magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< error_p >>
rect -103 0 -57 89
rect 57 0 103 89
rect 217 0 263 89
<< nmos >>
rect -28 0 28 89
rect 132 0 188 89
<< ndiff >>
rect -116 76 -28 89
rect -116 13 -103 76
rect -57 13 -28 76
rect -116 0 -28 13
rect 28 76 132 89
rect 28 13 57 76
rect 103 13 132 76
rect 28 0 132 13
rect 188 76 276 89
rect 188 13 217 76
rect 263 13 276 76
rect 188 0 276 13
<< ndiffc >>
rect -103 13 -57 76
rect 57 13 103 76
rect 217 13 263 76
<< polysilicon >>
rect -28 89 28 133
rect 132 89 188 133
rect -28 -44 28 0
rect 132 -44 188 0
<< metal1 >>
rect -103 76 -57 89
rect -103 0 -57 13
rect 57 76 103 89
rect 57 0 103 13
rect 217 76 263 89
rect 217 0 263 13
<< labels >>
flabel ndiffc 80 44 80 44 0 FreeSans 93 0 0 0 D
flabel ndiffc -68 44 -68 44 0 FreeSans 93 0 0 0 S
flabel ndiffc 227 44 227 44 0 FreeSans 93 0 0 0 S
<< end >>
