magic
tech gf180mcuD
magscale 1 10
timestamp 1765833244
<< nwell >>
rect -133 264 369 277
rect -133 -39 241 264
rect 242 -39 369 264
rect -133 -66 369 -39
<< polysilicon >>
rect -70 211 -15 245
rect 90 211 146 245
rect 251 211 307 245
rect -70 -34 -15 0
rect 90 -34 146 0
rect 251 -34 307 0
use pmos_5p04310591302013_3v256x8m81  pmos_5p04310591302013_3v256x8m81_0
timestamp 1765833244
transform 1 0 -14 0 1 0
box -230 -86 495 297
<< end >>
