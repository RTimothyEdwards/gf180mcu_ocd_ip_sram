magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< nwell >>
rect -426 -86 1422 1250
<< pmos >>
rect -252 0 -196 1164
rect -92 0 -36 1164
rect 69 0 125 1164
rect 229 0 285 1164
rect 390 0 446 1164
rect 550 0 606 1164
rect 711 0 767 1164
rect 871 0 927 1164
rect 1032 0 1088 1164
rect 1192 0 1248 1164
<< pdiff >>
rect -340 1151 -252 1164
rect -340 13 -327 1151
rect -281 13 -252 1151
rect -340 0 -252 13
rect -196 1151 -92 1164
rect -196 13 -167 1151
rect -121 13 -92 1151
rect -196 0 -92 13
rect -36 1151 69 1164
rect -36 13 -7 1151
rect 39 13 69 1151
rect -36 0 69 13
rect 125 1151 229 1164
rect 125 13 154 1151
rect 200 13 229 1151
rect 125 0 229 13
rect 285 1151 390 1164
rect 285 13 314 1151
rect 360 13 390 1151
rect 285 0 390 13
rect 446 1151 550 1164
rect 446 13 475 1151
rect 521 13 550 1151
rect 446 0 550 13
rect 606 1151 711 1164
rect 606 13 635 1151
rect 681 13 711 1151
rect 606 0 711 13
rect 767 1151 871 1164
rect 767 13 796 1151
rect 842 13 871 1151
rect 767 0 871 13
rect 927 1151 1032 1164
rect 927 13 956 1151
rect 1002 13 1032 1151
rect 927 0 1032 13
rect 1088 1151 1192 1164
rect 1088 13 1117 1151
rect 1163 13 1192 1151
rect 1088 0 1192 13
rect 1248 1151 1336 1164
rect 1248 13 1277 1151
rect 1323 13 1336 1151
rect 1248 0 1336 13
<< pdiffc >>
rect -327 13 -281 1151
rect -167 13 -121 1151
rect -7 13 39 1151
rect 154 13 200 1151
rect 314 13 360 1151
rect 475 13 521 1151
rect 635 13 681 1151
rect 796 13 842 1151
rect 956 13 1002 1151
rect 1117 13 1163 1151
rect 1277 13 1323 1151
<< polysilicon >>
rect -252 1164 -196 1208
rect -92 1164 -36 1208
rect 69 1164 125 1208
rect 229 1164 285 1208
rect 390 1164 446 1208
rect 550 1164 606 1208
rect 711 1164 767 1208
rect 871 1164 927 1208
rect 1032 1164 1088 1208
rect 1192 1164 1248 1208
rect -252 -44 -196 0
rect -92 -44 -36 0
rect 69 -44 125 0
rect 229 -44 285 0
rect 390 -44 446 0
rect 550 -44 606 0
rect 711 -44 767 0
rect 871 -44 927 0
rect 1032 -44 1088 0
rect 1192 -44 1248 0
<< metal1 >>
rect -327 1151 -281 1164
rect -327 0 -281 13
rect -167 1151 -121 1164
rect -167 0 -121 13
rect -7 1151 39 1164
rect -7 0 39 13
rect 154 1151 200 1164
rect 154 0 200 13
rect 314 1151 360 1164
rect 314 0 360 13
rect 475 1151 521 1164
rect 475 0 521 13
rect 635 1151 681 1164
rect 635 0 681 13
rect 796 1151 842 1164
rect 796 0 842 13
rect 956 1151 1002 1164
rect 956 0 1002 13
rect 1117 1151 1163 1164
rect 1117 0 1163 13
rect 1277 1151 1323 1164
rect 1277 0 1323 13
<< labels >>
flabel pdiffc 498 582 498 582 0 FreeSans 186 0 0 0 D
flabel pdiffc 349 582 349 582 0 FreeSans 186 0 0 0 S
flabel pdiffc 189 582 189 582 0 FreeSans 186 0 0 0 D
flabel pdiffc 28 582 28 582 0 FreeSans 186 0 0 0 S
flabel pdiffc -132 582 -132 582 0 FreeSans 186 0 0 0 D
flabel pdiffc -292 582 -292 582 0 FreeSans 186 0 0 0 S
flabel pdiffc 646 582 646 582 0 FreeSans 186 0 0 0 S
flabel pdiffc 807 582 807 582 0 FreeSans 186 0 0 0 D
flabel pdiffc 1128 582 1128 582 0 FreeSans 186 0 0 0 D
flabel pdiffc 967 582 967 582 0 FreeSans 186 0 0 0 S
flabel pdiffc 1288 582 1288 582 0 FreeSans 186 0 0 0 S
<< end >>
