magic
tech gf180mcuD
magscale 1 10
timestamp 1765833452
<< nwell >>
rect 4122 8232 9678 11499
rect 4701 5227 5502 5510
rect 4559 5188 5502 5227
rect 4545 5029 5502 5188
rect 379 4708 3801 4985
rect 379 4436 3957 4708
rect 3360 4193 3957 4436
rect 4351 4196 5502 5029
rect 7086 3606 7356 6533
rect 8225 3175 8240 5463
rect 9124 3272 9137 5463
rect -51 1571 6079 2400
rect 5543 596 6079 1571
rect 4995 -699 6079 596
<< nmos >>
rect 6672 183 6728 2300
rect 6832 183 6888 2300
rect 6992 183 7048 2300
rect 8414 2243 8470 2666
rect 8574 2243 8630 2666
rect 8734 2243 8790 2666
rect 8894 2243 8950 2666
rect 7515 338 7571 2031
rect 7675 338 7731 2031
rect 7835 338 7891 2031
rect 7995 338 8051 2031
<< pmos >>
rect 3550 4291 3606 4504
rect 3710 4291 3766 4504
<< ndiff >>
rect 6584 2287 6672 2300
rect 6584 208 6597 2287
rect 6643 208 6672 2287
rect 6584 183 6672 208
rect 6728 183 6832 2300
rect 6888 183 6992 2300
rect 7048 2287 7148 2300
rect 7048 208 7079 2287
rect 7125 208 7148 2287
rect 8323 2652 8414 2666
rect 8323 2338 8338 2652
rect 8385 2338 8414 2652
rect 8323 2243 8414 2338
rect 8470 2243 8574 2666
rect 8630 2652 8734 2666
rect 8630 2338 8659 2652
rect 8705 2338 8734 2652
rect 8630 2243 8734 2338
rect 8790 2243 8894 2666
rect 8950 2652 9044 2666
rect 8950 2338 8979 2652
rect 9025 2338 9044 2652
rect 8950 2243 9044 2338
rect 7424 2018 7515 2031
rect 7424 443 7438 2018
rect 7484 443 7515 2018
rect 7424 338 7515 443
rect 7571 338 7675 2031
rect 7731 2018 7835 2031
rect 7731 443 7760 2018
rect 7806 443 7835 2018
rect 7731 338 7835 443
rect 7891 338 7995 2031
rect 8051 2018 8144 2031
rect 8051 443 8080 2018
rect 8126 443 8144 2018
rect 8051 338 8144 443
rect 7048 183 7148 208
<< pdiff >>
rect 3455 4491 3550 4504
rect 3455 4317 3475 4491
rect 3521 4317 3550 4491
rect 3455 4291 3550 4317
rect 3606 4291 3710 4504
rect 3766 4490 3861 4504
rect 3766 4317 3795 4490
rect 3841 4317 3861 4490
rect 3766 4291 3861 4317
<< ndiffc >>
rect 6597 208 6643 2287
rect 7079 208 7125 2287
rect 8338 2338 8385 2652
rect 8659 2338 8705 2652
rect 8979 2338 9025 2652
rect 7438 443 7484 2018
rect 7760 443 7806 2018
rect 8080 443 8126 2018
<< pdiffc >>
rect 3475 4317 3521 4491
rect 3795 4317 3841 4490
<< psubdiff >>
rect 5593 8046 9620 8123
rect 5593 7858 5812 8046
rect 4437 4001 4531 4036
rect 4437 3840 4461 4001
rect 4507 3840 4531 4001
rect 4437 3500 4531 3840
<< nsubdiff >>
rect 4195 11398 9605 11423
rect 4195 11351 4327 11398
rect 9464 11351 9605 11398
rect 4195 11326 9605 11351
rect 4195 11271 4289 11326
rect 4195 8368 4219 11271
rect 4265 9212 4289 11271
rect 9511 11271 9605 11326
rect 4265 8404 6064 9212
rect 9511 8404 9535 11271
rect 4265 8379 9535 8404
rect 4265 8368 4327 8379
rect 4195 8333 4327 8368
rect 9464 8368 9535 8379
rect 9581 8368 9605 11271
rect 9464 8333 9605 8368
rect 4195 8308 9605 8333
rect 4437 4885 4531 4931
rect 4437 4455 4461 4885
rect 4507 4455 4531 4885
rect 4437 4349 4531 4455
<< psubdiffcont >>
rect 4461 3840 4507 4001
<< nsubdiffcont >>
rect 4327 11351 9464 11398
rect 4219 8368 4265 11271
rect 4327 8333 9464 8379
rect 9535 8368 9581 11271
rect 4461 4455 4507 4885
<< polysilicon >>
rect 4483 9315 4539 9393
rect 4643 9315 4699 9393
rect 4804 9315 4860 9393
rect 4964 9315 5020 9393
rect 5125 9315 5181 9393
rect 5285 9315 5341 9393
rect 5446 9315 5502 9393
rect 5606 9315 5662 9393
rect 5767 9315 5823 9393
rect 5927 9315 5983 9393
rect 6237 8562 6293 8845
rect 6397 8562 6453 8845
rect 6558 8562 6614 8845
rect 6718 8562 6774 8845
rect 6879 8562 6935 8845
rect 7039 8562 7095 8845
rect 7200 8562 7256 8845
rect 7360 8562 7416 8845
rect 7521 8562 7577 8845
rect 7681 8562 7737 8845
rect 7842 8562 7898 8845
rect 8002 8562 8058 8845
rect 8163 8562 8219 8845
rect 8323 8562 8379 8845
rect 8484 8562 8540 8845
rect 8645 8562 8701 8845
rect 8805 8562 8861 8845
rect 8966 8562 9022 8845
rect 9126 8562 9182 8845
rect 9287 8562 9343 8845
rect 6237 8487 9343 8562
rect 4695 7299 4751 7831
rect 4855 7299 4911 7831
rect 5016 7299 5072 7831
rect 5176 7299 5232 7831
rect 5337 7299 5393 7831
rect 6241 7614 6297 8024
rect 6401 7614 6457 8024
rect 6562 7614 6618 8024
rect 6722 7614 6778 8024
rect 6883 7614 6939 8024
rect 7043 7614 7099 8024
rect 7204 7614 7260 8024
rect 7364 7614 7420 8024
rect 7525 7614 7581 8024
rect 7685 7614 7741 8024
rect 7846 7614 7902 8024
rect 8006 7614 8062 8024
rect 8167 7614 8223 8024
rect 8327 7614 8383 8024
rect 8488 7614 8544 8024
rect 8649 7614 8705 8024
rect 8809 7614 8865 8024
rect 8970 7614 9026 8024
rect 9130 7614 9186 8024
rect 9291 7614 9347 8024
rect 3546 5289 3602 5519
rect 4893 5462 4949 5620
rect 5247 5572 5303 5617
rect 5247 5527 5537 5572
rect 4733 5217 4789 5272
rect 4893 5217 4949 5272
rect 4316 5175 4949 5217
rect 5247 5138 5303 5290
rect 3546 4986 3602 5005
rect 3546 4890 3763 4986
rect 3550 4504 3606 4656
rect 3710 4504 3766 4656
rect 5453 4884 5537 5527
rect 5247 4823 5537 4884
rect 5247 4713 5303 4823
rect 3550 3947 3606 4291
rect 3710 4099 3766 4291
rect 4733 4244 4789 4259
rect 4893 4244 4949 4259
rect 4733 4147 5077 4244
rect 5247 4158 5471 4201
rect 3710 4013 4106 4099
rect 3710 3947 3766 4013
rect 4733 4029 4789 4147
rect 4893 4029 4949 4147
rect 5247 4033 5303 4158
rect 3609 2282 3720 2633
rect 4364 2282 4475 2633
rect 4867 2303 4960 2657
rect 5320 2282 5376 2653
rect 5727 2523 5783 2750
rect 5727 2520 5905 2523
rect 5689 2425 5905 2520
rect 5689 2323 5745 2425
rect 5849 2324 5905 2425
rect 6672 2300 6728 3668
rect 6832 2300 6888 3668
rect 6992 2300 7048 3668
rect 7515 2031 7571 3221
rect 7675 2031 7731 3221
rect 7835 2031 7891 3221
rect 7995 2031 8051 3221
rect 8414 2666 8470 3221
rect 8574 2666 8630 3221
rect 8719 3108 8720 3167
rect 8734 2666 8790 3221
rect 8894 2666 8950 3221
rect 8414 2192 8470 2243
rect 8574 2192 8630 2243
rect 8734 2192 8790 2243
rect 8894 2192 8950 2243
rect 7515 288 7571 338
rect 7675 288 7731 338
rect 7835 288 7891 338
rect 7995 288 8051 338
rect 6672 133 6728 183
rect 6832 133 6888 183
rect 6992 133 7048 183
<< metal1 >>
rect 4202 11398 9599 11417
rect 4202 11351 4327 11398
rect 9464 11351 9599 11398
rect 4202 11333 9599 11351
rect 4202 11271 4489 11333
rect 4202 8368 4219 11271
rect 4265 9429 4489 11271
rect 4724 10237 4797 11333
rect 5045 10237 5118 11333
rect 5366 10237 5439 11333
rect 5687 10237 5760 11333
rect 6008 10237 6081 11333
rect 6159 10237 6232 11333
rect 6480 10237 6553 11333
rect 6801 10237 6874 11333
rect 7122 10237 7195 11333
rect 7443 10237 7516 11333
rect 7764 10237 7837 11333
rect 8085 10237 8158 11333
rect 8406 10237 8479 11333
rect 8727 10237 8800 11333
rect 9048 10237 9121 11333
rect 9310 11271 9599 11333
rect 4265 9198 4283 9429
rect 4265 8398 6051 9198
rect 9310 8603 9535 11271
rect 9517 8398 9535 8603
rect 4265 8379 9535 8398
rect 4265 8368 4327 8379
rect 4202 8333 4327 8368
rect 9464 8368 9535 8379
rect 9581 8368 9599 11271
rect 9464 8333 9599 8368
rect 4202 8314 9599 8333
rect 5607 7858 5798 8060
rect 4401 6926 4693 7717
rect 4402 6332 4693 6926
rect 9310 6892 9606 7864
rect 4402 6067 4483 6240
rect 248 5411 3004 6067
rect 3460 5980 3542 6064
rect 4401 5996 4483 6067
rect 5506 5983 5798 6067
rect 3461 5564 3542 5980
rect 4803 5800 5391 5873
rect 3618 5579 3699 5686
rect 3618 5450 3999 5579
rect 3461 4974 3542 5348
rect 3618 5042 3699 5450
rect 4646 5210 4727 5331
rect 4803 5283 4884 5800
rect 4960 5210 5041 5331
rect 4646 5139 5041 5210
rect 3460 4575 3542 4974
rect 3654 4895 3856 4980
rect 3461 4491 3542 4575
rect 3461 4317 3475 4491
rect 3521 4317 3542 4491
rect 3461 4298 3542 4317
rect 3775 4490 3856 4895
rect 3775 4317 3795 4490
rect 3841 4317 3856 4490
rect 3775 4093 3856 4317
rect 4443 4885 4727 4925
rect 4443 4455 4461 4885
rect 4507 4455 4727 4885
rect 4443 4301 4727 4455
rect 3461 4022 3856 4093
rect 3461 3783 3542 4022
rect 3617 3720 3699 3966
rect 3775 3786 3856 4022
rect 4443 4001 4727 4093
rect 4443 3840 4461 4001
rect 4507 3850 4727 4001
rect 4803 3879 4884 5044
rect 4960 4980 5041 5139
rect 4959 4866 5041 4980
rect 5163 4237 5244 5745
rect 5320 5329 5391 5800
rect 5298 5144 5511 5228
rect 4969 4153 5244 4237
rect 4507 3840 4524 3850
rect 3618 3615 3699 3720
rect 4443 3615 4524 3840
rect 4960 3615 5041 4029
rect 5163 3910 5244 4153
rect 5298 4001 5376 4781
rect 5455 4165 5511 5144
rect 5298 3917 6167 4001
rect 6263 3960 6672 6616
rect 6757 5521 6803 6334
rect 6904 5430 6986 6637
rect 7586 6588 7668 6637
rect 6591 3959 6672 3960
rect 5298 3787 5376 3917
rect 6087 3674 6167 3917
rect 7108 3705 7210 6435
rect 7587 5298 7668 6588
rect 7900 5315 7982 6637
rect 8486 5310 8567 6637
rect 8799 5305 8880 6637
rect 46 2933 5704 3615
rect 6086 3581 6167 3674
rect 5799 3417 6737 3501
rect 5799 2996 5880 3417
rect 3529 2682 3576 2933
rect 3770 2640 4101 2724
rect 4288 2640 4369 2933
rect 4020 2515 4101 2640
rect 4552 2515 4633 2742
rect 4793 2643 4847 2933
rect 5028 2515 5109 2742
rect 5243 2652 5324 2933
rect 5622 2764 5704 2933
rect 5404 2515 5451 2758
rect 5812 2574 5858 2808
rect 5772 2528 5858 2574
rect 4020 2431 4384 2515
rect 4552 2431 4890 2515
rect 5028 2431 5318 2515
rect 5404 2431 5702 2515
rect 3530 1918 3581 2285
rect 4020 2282 4101 2431
rect 4552 2293 4633 2431
rect 3750 2156 4101 2282
rect 3548 1733 3580 1918
rect 4281 1780 4363 2282
rect 4502 2197 4633 2293
rect 4788 1925 4869 2282
rect 5028 2198 5109 2431
rect 5243 1925 5324 2282
rect 5404 2193 5451 2431
rect 5419 2192 5451 2193
rect 4788 1908 5324 1925
rect 4788 1780 4869 1908
rect 4902 1634 5324 1908
rect 5602 1780 5684 2282
rect 5772 2192 5818 2528
rect 6214 2287 6672 3352
rect 7128 3287 7210 3705
rect 5916 1780 5997 2282
rect 4622 764 4670 860
rect 6214 208 6597 2287
rect 6643 208 6672 2287
rect 6214 -77 6672 208
rect 7061 3049 7210 3287
rect 8325 3201 8415 3298
rect 7508 3117 8415 3201
rect 8587 3094 9039 3178
rect 7061 2965 7880 3049
rect 7061 2287 7210 2965
rect 8158 2942 8959 3026
rect 7430 2822 7511 2872
rect 7061 208 7079 2287
rect 7125 208 7210 2287
rect 7061 189 7210 208
rect 7429 2018 7511 2822
rect 7429 443 7438 2018
rect 7484 443 7511 2018
rect 7743 2018 7825 2872
rect 7743 1561 7760 2018
rect 7429 139 7511 443
rect 7744 443 7760 1561
rect 7806 443 7825 2018
rect 7744 345 7825 443
rect 8057 2018 8138 2872
rect 8330 2822 8410 2872
rect 8057 443 8080 2018
rect 8126 443 8138 2018
rect 7430 25 7511 139
rect 7429 -46 7511 25
rect 8057 -77 8138 443
rect 8329 2652 8410 2822
rect 8329 2338 8338 2652
rect 8385 2338 8410 2652
rect 8329 139 8410 2338
rect 8642 2652 8724 2872
rect 8642 2338 8659 2652
rect 8705 2338 8724 2652
rect 8642 1561 8724 2338
rect 8956 2652 9523 2872
rect 8956 2338 8979 2652
rect 9025 2338 9523 2652
rect 8330 25 8410 139
rect 8329 -40 8410 25
rect 8956 -25 9523 2338
rect 6299 -588 9580 -268
<< metal2 >>
rect 4357 10234 9401 11394
rect 4559 9429 5903 10131
rect 4547 7774 5154 9363
rect 5313 8547 5734 9429
rect 6331 8751 9244 10063
rect 5313 7968 7811 8547
rect 4547 6234 4707 7774
rect 5313 7648 5734 7968
rect 8088 7897 9244 8751
rect 4766 7439 5734 7648
rect 5899 7511 9244 7897
rect 5899 6815 6103 7511
rect 6331 6815 6421 7511
rect 6645 6815 6735 7511
rect 6958 6815 7049 7511
rect 7272 6815 7362 7511
rect 7585 6815 7676 7511
rect 7899 6815 7989 7511
rect 8213 6815 8303 7511
rect 8526 6815 8617 7511
rect 8840 6815 8930 7511
rect 9153 6815 9244 7511
rect 5899 6548 9244 6815
rect 5899 6165 6103 6548
rect 3227 6061 6103 6165
rect 6743 6075 7148 6321
rect -196 5110 -102 5204
rect -195 -1217 -102 5110
rect 3299 4148 3393 6061
rect 3831 5518 3922 5996
rect 5455 5441 5545 5987
rect 3773 5269 5548 5366
rect 3773 4515 3866 5269
rect 4015 5110 4120 5202
rect 4016 3847 4120 5110
rect 4391 5004 4484 5189
rect 4391 4907 4872 5004
rect 5455 4981 5548 5269
rect 4862 4151 7070 4244
rect 4862 4150 4889 4151
rect 4016 3754 6911 3847
rect 4016 2519 4120 3754
rect 3892 2426 4120 2519
rect 6082 -177 6175 3674
rect 6821 3395 6911 3754
rect 6979 3398 7070 4151
rect 7224 -483 7315 6548
rect 8268 5988 9244 6548
rect 7743 3731 7825 5938
rect 7425 3408 8143 3731
rect 7744 3031 7825 3408
rect 8325 3266 9042 3817
rect 7744 2938 8327 3031
rect 7744 2872 7825 2938
rect 8643 2872 8724 3266
rect 7743 2639 7825 2872
rect 8642 2639 8724 2872
rect 9130 -483 9221 5988
<< metal3 >>
rect 1913 10180 9762 11398
rect 4190 6678 9762 7951
rect 4190 6657 7042 6678
rect 4547 6234 8138 6479
rect 8268 6007 10672 6557
rect 3761 5899 5618 5996
rect -144 5357 5653 5834
rect -223 5110 4186 5204
rect 5970 5001 9711 5908
rect 16 4390 9711 5001
rect 393 3720 9714 4246
rect 110 2853 6811 3496
rect 8817 3128 9056 3166
rect 8817 3099 9057 3128
rect 8976 3036 9057 3099
rect 8976 2970 9878 3036
rect 9812 2856 9878 2970
rect 110 2618 9648 2853
rect 9812 2790 11256 2856
rect 49 1585 6180 2328
rect 6456 1395 9648 2618
rect -313 1175 9648 1395
rect -651 976 9648 1175
rect -313 965 9648 976
rect -651 74 6010 272
rect 6456 126 9648 965
rect -12453 -607 12336 -289
rect -12453 -1055 11059 -810
rect -9940 -1218 11059 -1125
use M1_NACTIVE4310591302063_3v256x8m81  M1_NACTIVE4310591302063_3v256x8m81_0
timestamp 1763766357
transform 1 0 3915 0 1 1757
box -1288 -159 1288 159
use M1_NWELL01_3v256x8m81  M1_NWELL01_3v256x8m81_0
timestamp 1763766357
transform 1 0 1806 0 1 4709
box -1426 -273 1427 273
use M1_NWELL16_3v256x8m81  M1_NWELL16_3v256x8m81_0
timestamp 1763766357
transform -1 0 7798 0 -1 6630
box -1648 -158 1647 159
use M1_NWELL17_3v256x8m81  M1_NWELL17_3v256x8m81_0
timestamp 1763766357
transform 1 0 5235 0 1 8813
box -928 -501 928 501
use M1_NWELL_02_R90_3v256x8m81  M1_NWELL_02_R90_3v256x8m81_0
timestamp 1763766357
transform 0 -1 6358 1 0 5316
box -1473 -210 1473 209
use M1_NWELL_03_R90_3v256x8m81  M1_NWELL_03_R90_3v256x8m81_0
timestamp 1763766357
transform 0 -1 9347 1 0 5030
box -1758 -210 1759 210
use M1_PACTIVE01_3v256x8m81  M1_PACTIVE01_3v256x8m81_0
timestamp 1763766357
transform 1 0 2897 0 1 6025
box -2655 -56 2635 56
use M1_PACTIVE02_3v256x8m81  M1_PACTIVE02_3v256x8m81_0
timestamp 1763766357
transform -1 0 5051 0 -1 8018
box -662 -56 662 56
use M1_PACTIVE06_3v256x8m81  M1_PACTIVE06_3v256x8m81_0
timestamp 1763766357
transform 1 0 1806 0 1 4021
box -1326 -170 1327 170
use M1_PACTIVE4310591302068_3v256x8m81  M1_PACTIVE4310591302068_3v256x8m81_0
timestamp 1763766357
transform 1 0 2825 0 1 3271
box -2619 -239 2619 239
use M1_PACTIVE_01_R90_3v256x8m81  M1_PACTIVE_01_R90_3v256x8m81_0
timestamp 1763766357
transform 0 -1 4442 1 0 7104
box -965 -54 970 53
use M1_PACTIVE_02_R90_3v256x8m81  M1_PACTIVE_02_R90_3v256x8m81_0
timestamp 1764700137
transform 0 -1 9566 1 0 7529
box -627 -54 613 54
use M1_PACTIVE_03_R90_3v256x8m81  M1_PACTIVE_03_R90_3v256x8m81_0
timestamp 1763766357
transform 0 -1 5702 1 0 6939
box -970 -109 970 109
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_0
timestamp 1765833244
transform 1 0 5661 0 1 2473
box -67 -48 67 47
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_1
timestamp 1765833244
transform 1 0 5299 0 1 2473
box -67 -48 67 47
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_2
timestamp 1765833244
transform 1 0 4851 0 1 2473
box -67 -48 67 47
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_3
timestamp 1765833244
transform 1 0 5009 0 1 4195
box -67 -48 67 47
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_4
timestamp 1765833244
transform 1 0 5471 0 1 4207
box -67 -48 67 47
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_5
timestamp 1765833244
transform -1 0 3553 0 1 4200
box -67 -48 67 47
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_6
timestamp 1765833244
transform 1 0 4344 0 1 2473
box -67 -48 67 47
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_7
timestamp 1765833244
transform 1 0 3695 0 1 4938
box -67 -48 67 47
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_8
timestamp 1765833244
transform 1 0 5338 0 1 5186
box -67 -48 67 47
use M1_POLY2$$44754988_3v256x8m81  M1_POLY2$$44754988_3v256x8m81_0
timestamp 1765833244
transform -1 0 5496 0 1 5516
box -96 -124 67 124
use M1_POLY2$$46559276_3v256x8m81  M1_POLY2$$46559276_3v256x8m81_0
timestamp 1763766357
transform 1 0 3812 0 1 2473
box -123 -48 123 48
use M1_POLY2$$46559276_3v256x8m81  M1_POLY2$$46559276_3v256x8m81_1
timestamp 1763766357
transform 1 0 4439 0 1 5157
box -123 -48 123 48
use M1_POLY24310591302019_3v256x8m81  M1_POLY24310591302019_3v256x8m81_0
timestamp 1765833244
transform 1 0 6869 0 1 3517
box -36 -80 36 78
use M1_POLY24310591302019_3v256x8m81  M1_POLY24310591302019_3v256x8m81_1
timestamp 1765833244
transform 1 0 6713 0 1 3517
box -36 -80 36 78
use M1_POLY24310591302019_3v256x8m81  M1_POLY24310591302019_3v256x8m81_2
timestamp 1765833244
transform 1 0 7026 0 1 3517
box -36 -80 36 78
use M1_POLY24310591302030_3v256x8m81  M1_POLY24310591302030_3v256x8m81_0
timestamp 1765833244
transform 1 0 8687 0 1 3138
box -95 -36 95 36
use M1_POLY24310591302031_3v256x8m81  M1_POLY24310591302031_3v256x8m81_0
timestamp 1765833244
transform 1 0 8918 0 1 2985
box -36 -36 36 36
use M1_POLY24310591302031_3v256x8m81  M1_POLY24310591302031_3v256x8m81_1
timestamp 1765833244
transform 1 0 8448 0 1 2985
box -36 -36 36 36
use M1_POLY24310591302031_3v256x8m81  M1_POLY24310591302031_3v256x8m81_2
timestamp 1765833244
transform 1 0 8019 0 1 3159
box -36 -36 36 36
use M1_POLY24310591302031_3v256x8m81  M1_POLY24310591302031_3v256x8m81_3
timestamp 1765833244
transform 1 0 7550 0 1 3159
box -36 -36 36 36
use M1_POLY24310591302031_3v256x8m81  M1_POLY24310591302031_3v256x8m81_4
timestamp 1765833244
transform 1 0 4067 0 1 4051
box -36 -36 36 36
use M1_POLY24310591302033_3v256x8m81  M1_POLY24310591302033_3v256x8m81_0
timestamp 1765833244
transform 1 0 7783 0 1 3007
box -62 -36 62 36
use M1_POLY24310591302061_3v256x8m81  M1_POLY24310591302061_3v256x8m81_0
timestamp 1763766357
transform 1 0 7798 0 1 8526
box -1509 -36 1509 36
use M1_POLY24310591302062_3v256x8m81  M1_POLY24310591302062_3v256x8m81_0
timestamp 1764697366
transform 1 0 7776 0 1 7990
box -1550 -36 1550 36
use M1_POLY24310591302066_3v256x8m81  M1_POLY24310591302066_3v256x8m81_0
timestamp 1763766357
transform 1 0 5238 0 1 9351
box -720 -36 720 36
use M1_POLY24310591302067_3v256x8m81  M1_POLY24310591302067_3v256x8m81_0
timestamp 1763766357
transform 1 0 5048 0 1 7795
box -325 -36 325 36
use M1_PSUB$$48312364_3v256x8m81  M1_PSUB$$48312364_3v256x8m81_0
timestamp 1763766357
transform 1 0 7924 0 1 -25
box -1605 -58 1605 58
use M1_PSUB_02_R90_3v256x8m81  M1_PSUB_02_R90_3v256x8m81_0
timestamp 1763766357
transform 0 -1 6319 1 0 1631
box -1714 -111 1714 111
use M1_PSUB_03_3v256x8m81  M1_PSUB_03_3v256x8m81_0
timestamp 1763766357
transform -1 0 1626 0 1 5684
box -1383 -171 1383 172
use M1_PSUB_03_R90_3v256x8m81  M1_PSUB_03_R90_3v256x8m81_0
timestamp 1763766357
transform 0 -1 9418 1 0 1460
box -1543 -111 1542 111
use M2_M1$$34864172_3v256x8m81  M2_M1$$34864172_3v256x8m81_0
timestamp 1763766357
transform 1 0 8208 0 1 2984
box -119 -46 119 46
use M2_M1$$34864172_3v256x8m81  M2_M1$$34864172_3v256x8m81_1
timestamp 1763766357
transform 1 0 8935 0 1 3140
box -119 -46 119 46
use M2_M1$$34864172_3v256x8m81  M2_M1$$34864172_3v256x8m81_2
timestamp 1763766357
transform 1 0 3480 0 1 4195
box -119 -46 119 46
use M2_M1$$34864172_3v256x8m81  M2_M1$$34864172_3v256x8m81_3
timestamp 1763766357
transform 1 0 3845 0 1 2472
box -119 -46 119 46
use M2_M1$$34864172_R90_3v256x8m81  M2_M1$$34864172_R90_3v256x8m81_0
timestamp 1763766357
transform 0 -1 7025 1 0 3518
box -123 -45 123 45
use M2_M1$$34864172_R90_3v256x8m81  M2_M1$$34864172_R90_3v256x8m81_1
timestamp 1763766357
transform 0 -1 6867 1 0 3518
box -123 -45 123 45
use M2_M1$$34864172_R90_3v256x8m81  M2_M1$$34864172_R90_3v256x8m81_2
timestamp 1763766357
transform 0 -1 4844 1 0 4188
box -123 -45 123 45
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_0
timestamp 1765833244
transform 1 0 4488 0 1 4084
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_1
timestamp 1765833244
transform -1 0 3819 0 1 4616
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_2
timestamp 1765833244
transform -1 0 3658 0 1 3843
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_3
timestamp 1765833244
transform 1 0 6788 0 1 6198
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_4
timestamp 1765833244
transform 1 0 7103 0 1 6198
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_5
timestamp 1765833244
transform 1 0 5000 0 1 5612
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_6
timestamp 1765833244
transform 1 0 5499 0 1 5105
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_7
timestamp 1765833244
transform 1 0 5499 0 1 5563
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_8
timestamp 1765833244
transform 1 0 4844 0 1 4960
box -43 -122 43 122
use M2_M1$$43375660_R90_3v256x8m81  M2_M1$$43375660_R90_3v256x8m81_0
timestamp 1765833244
transform 0 -1 6128 1 0 3627
box -46 -119 46 119
use M2_M1$$43375660_R90_3v256x8m81  M2_M1$$43375660_R90_3v256x8m81_1
timestamp 1765833244
transform 0 -1 4426 1 0 5155
box -46 -119 46 119
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_0
timestamp 1763766357
transform 1 0 4448 0 1 10815
box -44 21 44 579
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_1
timestamp 1763766357
transform 1 0 4762 0 1 10815
box -44 21 44 579
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_2
timestamp 1763766357
transform 1 0 5075 0 1 10815
box -44 21 44 579
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_3
timestamp 1763766357
transform 1 0 5389 0 1 10815
box -44 21 44 579
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_4
timestamp 1763766357
transform 1 0 5702 0 1 10815
box -44 21 44 579
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_5
timestamp 1763766357
transform 1 0 6846 0 1 10815
box -44 21 44 579
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_6
timestamp 1763766357
transform 1 0 6533 0 1 10815
box -44 21 44 579
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_7
timestamp 1763766357
transform 1 0 6219 0 1 10815
box -44 21 44 579
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_8
timestamp 1763766357
transform 1 0 6016 0 1 10815
box -44 21 44 579
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_9
timestamp 1763766357
transform 1 0 8101 0 1 10815
box -44 21 44 579
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_10
timestamp 1763766357
transform 1 0 7787 0 1 10815
box -44 21 44 579
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_11
timestamp 1763766357
transform 1 0 7473 0 1 10815
box -44 21 44 579
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_12
timestamp 1763766357
transform 1 0 9355 0 1 10815
box -44 21 44 579
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_13
timestamp 1763766357
transform 1 0 9041 0 1 10815
box -44 21 44 579
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_14
timestamp 1763766357
transform 1 0 8728 0 1 10815
box -44 21 44 579
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_15
timestamp 1763766357
transform 1 0 8414 0 1 10815
box -44 21 44 579
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_16
timestamp 1763766357
transform 1 0 7160 0 1 10815
box -44 21 44 579
use M2_M1$$43377708_3v256x8m81  M2_M1$$43377708_3v256x8m81_0
timestamp 1763766357
transform 1 0 8885 0 1 7437
box -44 -427 44 427
use M2_M1$$43377708_3v256x8m81  M2_M1$$43377708_3v256x8m81_1
timestamp 1763766357
transform 1 0 7944 0 1 7437
box -44 -427 44 427
use M2_M1$$43377708_3v256x8m81  M2_M1$$43377708_3v256x8m81_2
timestamp 1763766357
transform 1 0 7630 0 1 7437
box -44 -427 44 427
use M2_M1$$43377708_3v256x8m81  M2_M1$$43377708_3v256x8m81_3
timestamp 1763766357
transform 1 0 7317 0 1 7437
box -44 -427 44 427
use M2_M1$$43377708_3v256x8m81  M2_M1$$43377708_3v256x8m81_4
timestamp 1763766357
transform 1 0 9198 0 1 7437
box -44 -427 44 427
use M2_M1$$43377708_3v256x8m81  M2_M1$$43377708_3v256x8m81_5
timestamp 1763766357
transform 1 0 8571 0 1 7437
box -44 -427 44 427
use M2_M1$$43377708_3v256x8m81  M2_M1$$43377708_3v256x8m81_6
timestamp 1763766357
transform 1 0 8257 0 1 7437
box -44 -427 44 427
use M2_M1$$43377708_3v256x8m81  M2_M1$$43377708_3v256x8m81_7
timestamp 1763766357
transform 1 0 7003 0 1 7437
box -44 -427 44 427
use M2_M1$$43377708_3v256x8m81  M2_M1$$43377708_3v256x8m81_8
timestamp 1763766357
transform 1 0 6376 0 1 7437
box -44 -427 44 427
use M2_M1$$43377708_3v256x8m81  M2_M1$$43377708_3v256x8m81_9
timestamp 1763766357
transform 1 0 6689 0 1 7437
box -44 -427 44 427
use M2_M1$$43378732_3v256x8m81  M2_M1$$43378732_3v256x8m81_0
timestamp 1763766357
transform 1 0 4603 0 1 9780
box -44 -351 44 351
use M2_M1$$43378732_3v256x8m81  M2_M1$$43378732_3v256x8m81_1
timestamp 1763766357
transform 1 0 5231 0 1 9780
box -44 -351 44 351
use M2_M1$$43378732_3v256x8m81  M2_M1$$43378732_3v256x8m81_2
timestamp 1763766357
transform 1 0 4917 0 1 9780
box -44 -351 44 351
use M2_M1$$43378732_3v256x8m81  M2_M1$$43378732_3v256x8m81_3
timestamp 1763766357
transform 1 0 5544 0 1 9780
box -44 -351 44 351
use M2_M1$$43378732_3v256x8m81  M2_M1$$43378732_3v256x8m81_4
timestamp 1763766357
transform 1 0 5858 0 1 9780
box -44 -351 44 351
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_0
timestamp 1763766357
transform 1 0 8997 0 1 3542
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_1
timestamp 1763766357
transform 1 0 8369 0 1 3542
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_2
timestamp 1763766357
transform 1 0 8683 0 1 3542
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_3
timestamp 1763766357
transform 1 0 9043 0 1 7168
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_4
timestamp 1763766357
transform 1 0 8102 0 1 7168
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_5
timestamp 1763766357
transform 1 0 8416 0 1 7168
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_6
timestamp 1763766357
transform 1 0 8729 0 1 7168
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_7
timestamp 1763766357
transform 1 0 7475 0 1 7168
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_8
timestamp 1763766357
transform 1 0 9566 0 1 7191
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_9
timestamp 1763766357
transform 1 0 7788 0 1 7168
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_10
timestamp 1763766357
transform 1 0 9355 0 1 7168
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_11
timestamp 1763766357
transform 1 0 4967 0 1 6936
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_12
timestamp 1763766357
transform 1 0 6848 0 1 7168
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_13
timestamp 1763766357
transform 1 0 6534 0 1 7168
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_14
timestamp 1763766357
transform 1 0 6220 0 1 7168
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_15
timestamp 1763766357
transform 1 0 5280 0 1 6936
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_16
timestamp 1763766357
transform 1 0 7161 0 1 7168
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_17
timestamp 1763766357
transform 1 0 5000 0 1 4705
box -44 -275 44 275
use M2_M1$$43380780_3v256x8m81  M2_M1$$43380780_3v256x8m81_0
timestamp 1763766357
transform 1 0 4488 0 1 4629
box -44 -198 44 198
use M2_M1$$43380780_3v256x8m81  M2_M1$$43380780_3v256x8m81_1
timestamp 1763766357
transform -1 0 3501 0 1 4774
box -44 -198 44 198
use M2_M1$$45013036_3v256x8m81  M2_M1$$45013036_3v256x8m81_0
timestamp 1765833244
transform 1 0 4844 0 1 9317
box -266 -46 266 46
use M2_M1$$45013036_3v256x8m81  M2_M1$$45013036_3v256x8m81_1
timestamp 1765833244
transform 1 0 4865 0 1 7821
box -266 -46 266 46
use M2_M1$$47500332_3v256x8m81  M2_M1$$47500332_3v256x8m81_0
timestamp 1763766357
transform 1 0 9398 0 1 5176
box -44 -432 44 732
use M2_M1$$47500332_3v256x8m81  M2_M1$$47500332_3v256x8m81_1
timestamp 1763766357
transform 1 0 8525 0 1 5176
box -44 -432 44 732
use M2_M1$$47500332_3v256x8m81  M2_M1$$47500332_3v256x8m81_2
timestamp 1763766357
transform 1 0 8838 0 1 5176
box -44 -432 44 732
use M2_M1$$47500332_3v256x8m81  M2_M1$$47500332_3v256x8m81_3
timestamp 1763766357
transform 1 0 6945 0 1 5173
box -44 -432 44 732
use M2_M1$$47500332_3v256x8m81  M2_M1$$47500332_3v256x8m81_4
timestamp 1763766357
transform 1 0 6631 0 1 5173
box -44 -432 44 732
use M2_M1$$47500332_3v256x8m81  M2_M1$$47500332_3v256x8m81_5
timestamp 1763766357
transform 1 0 7941 0 1 5166
box -44 -432 44 732
use M2_M1$$47500332_3v256x8m81  M2_M1$$47500332_3v256x8m81_6
timestamp 1763766357
transform 1 0 7627 0 1 5166
box -44 -432 44 732
use M2_M1$$47515692_3v256x8m81  M2_M1$$47515692_3v256x8m81_0
timestamp 1763766357
transform 1 0 4438 0 1 7429
box -44 -504 44 284
use M2_M1$$47515692_3v256x8m81  M2_M1$$47515692_3v256x8m81_1
timestamp 1763766357
transform 1 0 4810 0 1 7165
box -44 -504 44 284
use M2_M1$$47515692_3v256x8m81  M2_M1$$47515692_3v256x8m81_2
timestamp 1763766357
transform 1 0 5436 0 1 7165
box -44 -504 44 284
use M2_M1$$47515692_3v256x8m81  M2_M1$$47515692_3v256x8m81_3
timestamp 1763766357
transform 1 0 5123 0 1 7165
box -44 -504 44 284
use M2_M1$$48217132_3v256x8m81  M2_M1$$48217132_3v256x8m81_0
timestamp 1763766357
transform 1 0 7784 0 1 2216
box -44 -655 45 655
use M2_M1$$48217132_3v256x8m81  M2_M1$$48217132_3v256x8m81_1
timestamp 1763766357
transform 1 0 8683 0 1 2216
box -44 -655 45 655
use M2_M1$$48217132_3v256x8m81  M2_M1$$48217132_3v256x8m81_2
timestamp 1763766357
transform 1 0 7003 0 1 9407
box -44 -655 45 655
use M2_M1$$48217132_3v256x8m81  M2_M1$$48217132_3v256x8m81_3
timestamp 1763766357
transform 1 0 6689 0 1 9407
box -44 -655 45 655
use M2_M1$$48217132_3v256x8m81  M2_M1$$48217132_3v256x8m81_4
timestamp 1763766357
transform 1 0 6376 0 1 9407
box -44 -655 45 655
use M2_M1$$48217132_3v256x8m81  M2_M1$$48217132_3v256x8m81_5
timestamp 1763766357
transform 1 0 9198 0 1 9407
box -44 -655 45 655
use M2_M1$$48217132_3v256x8m81  M2_M1$$48217132_3v256x8m81_6
timestamp 1763766357
transform 1 0 8257 0 1 9407
box -44 -655 45 655
use M2_M1$$48217132_3v256x8m81  M2_M1$$48217132_3v256x8m81_7
timestamp 1763766357
transform 1 0 8571 0 1 9407
box -44 -655 45 655
use M2_M1$$48217132_3v256x8m81  M2_M1$$48217132_3v256x8m81_8
timestamp 1763766357
transform 1 0 8885 0 1 9407
box -44 -655 45 655
use M2_M1$$48217132_3v256x8m81  M2_M1$$48217132_3v256x8m81_9
timestamp 1763766357
transform 1 0 7317 0 1 9407
box -44 -655 45 655
use M2_M1$$48217132_3v256x8m81  M2_M1$$48217132_3v256x8m81_10
timestamp 1763766357
transform 1 0 7630 0 1 9407
box -44 -655 45 655
use M2_M1$$48217132_3v256x8m81  M2_M1$$48217132_3v256x8m81_11
timestamp 1763766357
transform 1 0 7944 0 1 9407
box -44 -655 45 655
use M2_M1$$48218156_3v256x8m81  M2_M1$$48218156_3v256x8m81_0
timestamp 1763766357
transform 1 0 7081 0 1 8500
box -709 -46 709 46
use M2_M1$$48218156_3v256x8m81  M2_M1$$48218156_3v256x8m81_1
timestamp 1763766357
transform 1 0 7081 0 1 8015
box -709 -46 709 46
use M2_M1$$48219180_3v256x8m81  M2_M1$$48219180_3v256x8m81_0
timestamp 1763766357
transform 1 0 6379 0 1 3043
box -119 -275 119 275
use M2_M1$$48220204_3v256x8m81  M2_M1$$48220204_3v256x8m81_0
timestamp 1763766357
transform 1 0 6376 0 1 5173
box -119 -732 119 732
use M2_M1$$48221228_3v256x8m81  M2_M1$$48221228_3v256x8m81_0
timestamp 1763766357
transform 1 0 9478 0 1 1480
box -44 -1341 45 1341
use M2_M1$$48221228_3v256x8m81  M2_M1$$48221228_3v256x8m81_1
timestamp 1763766357
transform 1 0 8098 0 1 1480
box -44 -1341 45 1341
use M2_M1$$48221228_3v256x8m81  M2_M1$$48221228_3v256x8m81_2
timestamp 1763766357
transform 1 0 8369 0 1 1480
box -44 -1341 45 1341
use M2_M1$$48221228_3v256x8m81  M2_M1$$48221228_3v256x8m81_3
timestamp 1763766357
transform 1 0 8997 0 1 1480
box -44 -1341 45 1341
use M2_M1$$48221228_3v256x8m81  M2_M1$$48221228_3v256x8m81_4
timestamp 1763766357
transform 1 0 7471 0 1 1480
box -44 -1341 45 1341
use M2_M1$$48222252_3v256x8m81  M2_M1$$48222252_3v256x8m81_0
timestamp 1763766357
transform 1 0 8098 0 1 4902
box -45 -1493 45 1493
use M2_M1$$48222252_3v256x8m81  M2_M1$$48222252_3v256x8m81_1
timestamp 1763766357
transform 1 0 7471 0 1 4902
box -45 -1493 45 1493
use M2_M1$$48222252_3v256x8m81  M2_M1$$48222252_3v256x8m81_2
timestamp 1763766357
transform 1 0 7784 0 1 4902
box -45 -1493 45 1493
use M2_M1$$48224300_3v256x8m81  M2_M1$$48224300_3v256x8m81_0
timestamp 1763766357
transform 1 0 5704 0 1 7009
box -118 -351 119 351
use M2_M1$$48316460_3v256x8m81  M2_M1$$48316460_3v256x8m81_0
timestamp 1763766357
transform 1 0 6636 0 1 1772
box -45 -1570 45 1570
use M2_M1$$168351788_3v256x8m81  M2_M1$$168351788_3v256x8m81_0
timestamp 1763766357
transform 1 0 4070 0 1 3970
box -45 -123 45 123
use M2_M1$$170061868_3v256x8m81  M2_M1$$170061868_3v256x8m81_0
timestamp 1763766357
transform 1 0 1967 0 1 3208
box -1815 -275 1815 275
use M2_M1$$170063916_3v256x8m81  M2_M1$$170063916_3v256x8m81_0
timestamp 1763766357
transform -1 0 1592 0 1 5609
box -1299 -198 1299 198
use M2_M1$$170064940_3v256x8m81  M2_M1$$170064940_3v256x8m81_0
timestamp 1763766357
transform -1 0 1792 0 1 4019
box -1299 -123 1299 123
use M2_M1$$170064940_3v256x8m81  M2_M1$$170064940_3v256x8m81_1
timestamp 1763766357
transform -1 0 1792 0 1 4708
box -1299 -123 1299 123
use M2_M1$$199746604_3v256x8m81  M2_M1$$199746604_3v256x8m81_0
timestamp 1763766357
transform 1 0 7269 0 1 -428
box -119 -123 119 123
use M2_M1$$199746604_3v256x8m81  M2_M1$$199746604_3v256x8m81_1
timestamp 1763766357
transform 1 0 9175 0 1 -428
box -119 -123 119 123
use M2_M1_01_R270_3v256x8m81  M2_M1_01_R270_3v256x8m81_0
timestamp 1763766357
transform 0 -1 3880 -1 0 5520
box -46 -119 46 119
use M2_M14310591302025_3v256x8m81  M2_M14310591302025_3v256x8m81_0
timestamp 1765833244
transform 1 0 5643 0 1 2016
box -34 -85 34 135
use M2_M14310591302025_3v256x8m81  M2_M14310591302025_3v256x8m81_1
timestamp 1765833244
transform 1 0 5957 0 1 2016
box -34 -85 34 135
use M2_M14310591302065_3v256x8m81  M2_M14310591302065_3v256x8m81_0
timestamp 1763766357
transform 1 0 3542 0 1 1754
box -1782 -165 1782 165
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_0
timestamp 1763766357
transform 1 0 4488 0 1 4084
box -44 -123 44 123
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_1
timestamp 1763766357
transform -1 0 3658 0 1 3843
box -44 -123 44 123
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_2
timestamp 1763766357
transform 1 0 8098 0 1 6357
box -44 -123 44 123
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_3
timestamp 1763766357
transform 1 0 7784 0 1 6357
box -44 -123 44 123
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_4
timestamp 1763766357
transform 1 0 7469 0 1 6357
box -44 -123 44 123
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_5
timestamp 1763766357
transform 1 0 5000 0 1 5612
box -44 -123 44 123
use M3_M2$$43368492_R270_3v256x8m81  M3_M2$$43368492_R270_3v256x8m81_0
timestamp 1763766357
transform 0 -1 3880 -1 0 5949
box -46 -119 46 119
use M3_M2$$43368492_R270_3v256x8m81  M3_M2$$43368492_R270_3v256x8m81_1
timestamp 1763766357
transform 0 -1 5499 -1 0 5949
box -46 -119 46 119
use M3_M2$$43371564_3v256x8m81  M3_M2$$43371564_3v256x8m81_0
timestamp 1765833244
transform 1 0 8935 0 1 3140
box -119 -46 119 46
use M3_M2$$43371564_3v256x8m81  M3_M2$$43371564_3v256x8m81_1
timestamp 1765833244
transform 1 0 -104 0 1 5157
box -119 -46 119 46
use M3_M2$$43371564_3v256x8m81  M3_M2$$43371564_3v256x8m81_2
timestamp 1765833244
transform 1 0 3346 0 1 6112
box -119 -46 119 46
use M3_M2$$43371564_3v256x8m81  M3_M2$$43371564_3v256x8m81_3
timestamp 1765833244
transform 1 0 4067 0 1 5157
box -119 -46 119 46
use M3_M2$$45008940_3v256x8m81  M3_M2$$45008940_3v256x8m81_0
timestamp 1765833244
transform 1 0 4702 0 1 6357
box -119 -123 119 123
use M3_M2$$47108140_3v256x8m81  M3_M2$$47108140_3v256x8m81_0
timestamp 1763766357
transform 1 0 4488 0 1 4629
box -45 -198 45 198
use M3_M2$$47108140_3v256x8m81  M3_M2$$47108140_3v256x8m81_1
timestamp 1763766357
transform -1 0 3501 0 1 4774
box -45 -198 45 198
use M3_M2$$47115308_3v256x8m81  M3_M2$$47115308_3v256x8m81_0
timestamp 1763766357
transform 1 0 6379 0 1 3043
box -119 -275 119 275
use M3_M2$$47332396_3v256x8m81  M3_M2$$47332396_3v256x8m81_0
timestamp 1763766357
transform 1 0 4438 0 1 7429
box -45 -504 45 504
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_0
timestamp 1763766357
transform 1 0 9355 0 1 7168
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_1
timestamp 1763766357
transform 1 0 7788 0 1 7168
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_2
timestamp 1763766357
transform 1 0 7475 0 1 7168
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_3
timestamp 1763766357
transform 1 0 8729 0 1 7168
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_4
timestamp 1763766357
transform 1 0 9566 0 1 7191
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_5
timestamp 1763766357
transform 1 0 8416 0 1 7168
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_6
timestamp 1763766357
transform 1 0 8102 0 1 7168
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_7
timestamp 1763766357
transform 1 0 9043 0 1 7168
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_8
timestamp 1763766357
transform 1 0 5280 0 1 6936
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_9
timestamp 1763766357
transform 1 0 6220 0 1 7168
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_10
timestamp 1763766357
transform 1 0 6534 0 1 7168
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_11
timestamp 1763766357
transform 1 0 6848 0 1 7168
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_12
timestamp 1763766357
transform 1 0 4967 0 1 6936
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_13
timestamp 1763766357
transform 1 0 7161 0 1 7168
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_14
timestamp 1763766357
transform 1 0 5000 0 1 4705
box -84 -185 84 275
use M3_M2$$47644716_3v256x8m81  M3_M2$$47644716_3v256x8m81_0
timestamp 1763766357
transform 1 0 8525 0 1 5176
box -45 -432 45 732
use M3_M2$$47644716_3v256x8m81  M3_M2$$47644716_3v256x8m81_1
timestamp 1763766357
transform 1 0 8838 0 1 5176
box -45 -432 45 732
use M3_M2$$47644716_3v256x8m81  M3_M2$$47644716_3v256x8m81_2
timestamp 1763766357
transform 1 0 6945 0 1 5173
box -45 -432 45 732
use M3_M2$$47644716_3v256x8m81  M3_M2$$47644716_3v256x8m81_3
timestamp 1763766357
transform 1 0 6631 0 1 5173
box -45 -432 45 732
use M3_M2$$47644716_3v256x8m81  M3_M2$$47644716_3v256x8m81_4
timestamp 1763766357
transform 1 0 7941 0 1 5166
box -45 -432 45 732
use M3_M2$$47644716_3v256x8m81  M3_M2$$47644716_3v256x8m81_5
timestamp 1763766357
transform 1 0 7627 0 1 5166
box -45 -432 45 732
use M3_M2$$47644716_3v256x8m81  M3_M2$$47644716_3v256x8m81_6
timestamp 1763766357
transform 1 0 9398 0 1 5176
box -45 -432 45 732
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_0
timestamp 1763766357
transform 1 0 4448 0 1 10815
box -45 -579 45 579
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_1
timestamp 1763766357
transform 1 0 5075 0 1 10815
box -45 -579 45 579
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_2
timestamp 1763766357
transform 1 0 5389 0 1 10815
box -45 -579 45 579
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_3
timestamp 1763766357
transform 1 0 5702 0 1 10815
box -45 -579 45 579
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_4
timestamp 1763766357
transform 1 0 6219 0 1 10815
box -45 -579 45 579
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_5
timestamp 1763766357
transform 1 0 6846 0 1 10815
box -45 -579 45 579
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_6
timestamp 1763766357
transform 1 0 6533 0 1 10815
box -45 -579 45 579
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_7
timestamp 1763766357
transform 1 0 6016 0 1 10815
box -45 -579 45 579
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_8
timestamp 1763766357
transform 1 0 4762 0 1 10815
box -45 -579 45 579
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_9
timestamp 1763766357
transform 1 0 7473 0 1 10815
box -45 -579 45 579
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_10
timestamp 1763766357
transform 1 0 9355 0 1 10815
box -45 -579 45 579
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_11
timestamp 1763766357
transform 1 0 9041 0 1 10815
box -45 -579 45 579
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_12
timestamp 1763766357
transform 1 0 8728 0 1 10815
box -45 -579 45 579
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_13
timestamp 1763766357
transform 1 0 8414 0 1 10815
box -45 -579 45 579
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_14
timestamp 1763766357
transform 1 0 8101 0 1 10815
box -45 -579 45 579
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_15
timestamp 1763766357
transform 1 0 7787 0 1 10815
box -45 -579 45 579
use M3_M2$$47645740_3v256x8m81  M3_M2$$47645740_3v256x8m81_16
timestamp 1763766357
transform 1 0 7160 0 1 10815
box -45 -579 45 579
use M3_M2$$48066604_3v256x8m81  M3_M2$$48066604_3v256x8m81_0
timestamp 1763766357
transform 1 0 8755 0 1 6282
box -487 -275 487 275
use M3_M2$$48227372_3v256x8m81  M3_M2$$48227372_3v256x8m81_0
timestamp 1763766357
transform 1 0 6636 0 1 1772
box -45 -1570 45 1570
use M3_M2$$48228396_3v256x8m81  M3_M2$$48228396_3v256x8m81_0
timestamp 1763766357
transform 1 0 6376 0 1 5173
box -119 -732 119 732
use M3_M2$$48229420_3v256x8m81  M3_M2$$48229420_3v256x8m81_0
timestamp 1763766357
transform 1 0 8098 0 1 1480
box -45 -1341 45 1341
use M3_M2$$48229420_3v256x8m81  M3_M2$$48229420_3v256x8m81_1
timestamp 1763766357
transform 1 0 8369 0 1 1480
box -45 -1341 45 1341
use M3_M2$$48229420_3v256x8m81  M3_M2$$48229420_3v256x8m81_2
timestamp 1763766357
transform 1 0 8997 0 1 1480
box -45 -1341 45 1341
use M3_M2$$48229420_3v256x8m81  M3_M2$$48229420_3v256x8m81_3
timestamp 1763766357
transform 1 0 7471 0 1 1480
box -45 -1341 45 1341
use M3_M2$$48229420_3v256x8m81  M3_M2$$48229420_3v256x8m81_4
timestamp 1763766357
transform 1 0 9478 0 1 1480
box -45 -1341 45 1341
use M3_M2$$48231468_3v256x8m81  M3_M2$$48231468_3v256x8m81_0
timestamp 1763766357
transform 1 0 5704 0 1 7009
box -119 -351 119 351
use M3_M2$$169753644_3v256x8m81  M3_M2$$169753644_3v256x8m81_0
timestamp 1763766357
transform 1 0 1967 0 1 3208
box -1815 -275 1815 275
use M3_M2$$169755692_3v256x8m81  M3_M2$$169755692_3v256x8m81_0
timestamp 1763766357
transform -1 0 1592 0 1 5609
box -1299 -198 1299 198
use M3_M2$$169756716_3v256x8m81  M3_M2$$169756716_3v256x8m81_0
timestamp 1763766357
transform -1 0 1792 0 1 4708
box -1299 -123 1299 123
use M3_M2$$169756716_3v256x8m81  M3_M2$$169756716_3v256x8m81_1
timestamp 1763766357
transform -1 0 1792 0 1 4019
box -1299 -123 1299 123
use M3_M2$$201255980_3v256x8m81  M3_M2$$201255980_3v256x8m81_0
timestamp 1763766357
transform 1 0 -149 0 1 -1171
box -119 -46 119 46
use M3_M24310591302026_3v256x8m81  M3_M24310591302026_3v256x8m81_0
timestamp 1765833244
transform 1 0 5643 0 1 2016
box -35 -135 35 135
use M3_M24310591302026_3v256x8m81  M3_M24310591302026_3v256x8m81_1
timestamp 1765833244
transform 1 0 5957 0 1 2016
box -35 -135 35 135
use M3_M24310591302064_3v256x8m81  M3_M24310591302064_3v256x8m81_0
timestamp 1763766357
transform 1 0 3542 0 1 1754
box -1782 -165 1782 165
use nmos_1p2$$46551084_3v256x8m81  nmos_1p2$$46551084_3v256x8m81_0
timestamp 1765833452
transform 1 0 5261 0 1 3781
box -102 -44 130 255
use nmos_1p2$$46563372_3v256x8m81  nmos_1p2$$46563372_3v256x8m81_0
timestamp 1765833452
transform 1 0 3560 0 1 5558
box -102 -44 130 133
use nmos_1p2$$46563372_3v256x8m81  nmos_1p2$$46563372_3v256x8m81_1
timestamp 1765833452
transform 1 0 4907 0 -1 5749
box -102 -44 130 133
use nmos_1p2$$46563372_3v256x8m81  nmos_1p2$$46563372_3v256x8m81_2
timestamp 1765833452
transform 1 0 5261 0 -1 5749
box -102 -44 130 133
use nmos_1p2$$47342636_3v256x8m81  nmos_1p2$$47342636_3v256x8m81_0
timestamp 1763766357
transform 1 0 3724 0 1 3781
box -102 -44 130 170
use nmos_1p2$$47342636_3v256x8m81  nmos_1p2$$47342636_3v256x8m81_1
timestamp 1763766357
transform 1 0 3564 0 1 3781
box -102 -44 130 170
use nmos_1p2$$48302124_3v256x8m81  nmos_1p2$$48302124_3v256x8m81_0
timestamp 1763766357
transform 1 0 5741 0 -1 3075
box -102 -44 130 325
use nmos_1p2$$48306220_3v256x8m81  nmos_1p2$$48306220_3v256x8m81_0
timestamp 1763766357
transform 1 0 4821 0 1 6327
box -214 -44 660 975
use nmos_1p2$$48308268_3v256x8m81  nmos_1p2$$48308268_3v256x8m81_0
timestamp 1763766357
transform 1 0 6787 0 1 6887
box -634 -44 2648 731
use nmos_1p2$$48629804_3v256x8m81  nmos_1p2$$48629804_3v256x8m81_0
timestamp 1765833452
transform 1 0 4775 0 1 3781
box -130 -44 262 255
use nmos_5p04310591302083_3v256x8m81  nmos_5p04310591302083_3v256x8m81_0
timestamp 1763766357
transform 1 0 5320 0 -1 2758
box -92 -44 148 114
use nmos_5p04310591302090_3v256x8m81  nmos_5p04310591302090_3v256x8m81_0
timestamp 1763766357
transform 1 0 4867 0 -1 2727
box -92 -44 185 100
use nmos_5p04310591302093_3v256x8m81  nmos_5p04310591302093_3v256x8m81_0
timestamp 1763766357
transform 1 0 3609 0 -1 2724
box -92 -44 204 100
use nmos_5p04310591302093_3v256x8m81  nmos_5p04310591302093_3v256x8m81_1
timestamp 1763766357
transform 1 0 4364 0 -1 2724
box -92 -44 204 100
use pmos_1p2$$46273580_3v256x8m81  pmos_1p2$$46273580_3v256x8m81_0
timestamp 1765833244
transform 1 0 4775 0 -1 5419
box -216 -86 348 192
use pmos_1p2$$46285868_3v256x8m81  pmos_1p2$$46285868_3v256x8m81_0
timestamp 1765833452
transform 1 0 3560 0 1 5036
box -188 -86 216 297
use pmos_1p2$$46285868_3v256x8m81  pmos_1p2$$46285868_3v256x8m81_1
timestamp 1765833452
transform 1 0 5261 0 1 4463
box -188 -86 216 297
use pmos_1p2$$47330348_3v256x8m81  pmos_1p2$$47330348_3v256x8m81_0
timestamp 1765833452
transform 1 0 5261 0 -1 5419
box -188 -86 216 175
use pmos_1p2$$47815724_3v256x8m81  pmos_1p2$$47815724_3v256x8m81_0
timestamp 1763766357
transform 1 0 8748 0 1 3261
box -188 -86 216 2202
use pmos_1p2$$47815724_3v256x8m81  pmos_1p2$$47815724_3v256x8m81_1
timestamp 1763766357
transform 1 0 8908 0 1 3261
box -188 -86 216 2202
use pmos_1p2$$47815724_3v256x8m81  pmos_1p2$$47815724_3v256x8m81_2
timestamp 1763766357
transform 1 0 8588 0 1 3261
box -188 -86 216 2202
use pmos_1p2$$47815724_3v256x8m81  pmos_1p2$$47815724_3v256x8m81_3
timestamp 1763766357
transform 1 0 8428 0 1 3261
box -188 -86 216 2202
use pmos_1p2$$47815724_3v256x8m81  pmos_1p2$$47815724_3v256x8m81_4
timestamp 1763766357
transform 1 0 8009 0 1 3261
box -188 -86 216 2202
use pmos_1p2$$47815724_3v256x8m81  pmos_1p2$$47815724_3v256x8m81_5
timestamp 1763766357
transform 1 0 7689 0 1 3261
box -188 -86 216 2202
use pmos_1p2$$47815724_3v256x8m81  pmos_1p2$$47815724_3v256x8m81_6
timestamp 1763766357
transform 1 0 7529 0 1 3261
box -188 -86 216 2202
use pmos_1p2$$47815724_3v256x8m81  pmos_1p2$$47815724_3v256x8m81_7
timestamp 1763766357
transform 1 0 7849 0 1 3261
box -188 -86 216 2202
use pmos_1p2$$48623660_3v256x8m81  pmos_1p2$$48623660_3v256x8m81_0
timestamp 1763766357
transform 1 0 5731 0 -1 2282
box -216 -86 348 437
use pmos_1p2$$48624684_3v256x8m81  pmos_1p2$$48624684_3v256x8m81_0
timestamp 1763766357
transform 1 0 7006 0 1 3705
box -188 -86 216 1906
use pmos_1p2$$48624684_3v256x8m81  pmos_1p2$$48624684_3v256x8m81_1
timestamp 1763766357
transform 1 0 6686 0 1 3705
box -188 -86 216 1906
use pmos_1p2$$48624684_3v256x8m81  pmos_1p2$$48624684_3v256x8m81_2
timestamp 1763766357
transform 1 0 6846 0 1 3705
box -188 -86 216 1906
use pmos_5p04310591302051_3v256x8m81  pmos_5p04310591302051_3v256x8m81_0
timestamp 1765833244
transform 1 0 4761 0 1 4295
box -202 -86 362 615
use pmos_5p04310591302074_3v256x8m81  pmos_5p04310591302074_3v256x8m81_0
timestamp 1763766357
transform 1 0 3609 0 -1 2282
box -174 -86 286 170
use pmos_5p04310591302074_3v256x8m81  pmos_5p04310591302074_3v256x8m81_1
timestamp 1763766357
transform 1 0 4364 0 -1 2282
box -174 -86 286 170
use pmos_5p04310591302088_3v256x8m81  pmos_5p04310591302088_3v256x8m81_0
timestamp 1763766357
transform 1 0 4735 0 1 9432
box -426 -86 1422 1250
use pmos_5p04310591302089_3v256x8m81  pmos_5p04310591302089_3v256x8m81_0
timestamp 1763766357
transform 1 0 6785 0 1 8878
box -722 -86 2732 1800
use pmos_5p04310591302092_3v256x8m81  pmos_5p04310591302092_3v256x8m81_0
timestamp 1763766357
transform 1 0 4867 0 -1 2282
box -174 -86 267 170
use pmos_5p04310591302094_3v256x8m81  pmos_5p04310591302094_3v256x8m81_0
timestamp 1763766357
transform 1 0 5320 0 -1 2282
box -174 -86 230 262
use wen_v2_3v256x8m81  wen_v2_3v256x8m81_0
timestamp 1765833452
transform 1 0 -11 0 1 -1312
box -30 -62 5184 2488
<< labels >>
flabel metal3 s 592 4041 592 4041 0 FreeSans 700 0 0 0 VSS
port 1 nsew
flabel metal3 s 224 2807 224 2807 0 FreeSans 700 0 0 0 VSS
port 1 nsew
flabel metal3 s 300 4674 300 4674 0 FreeSans 700 0 0 0 VDD
port 2 nsew
flabel metal3 s 592 5635 592 5635 0 FreeSans 700 0 0 0 VSS
port 1 nsew
flabel metal3 s 4489 7046 4489 7046 0 FreeSans 700 0 0 0 VSS
port 1 nsew
flabel metal3 s 240 1719 240 1719 0 FreeSans 700 0 0 0 VDD
port 2 nsew
flabel metal3 s 4489 10789 4489 10789 0 FreeSans 700 0 0 0 VDD
port 2 nsew
flabel metal3 s 1528 637 1528 637 0 FreeSans 700 0 0 0 IGWEN
port 4 nsew
rlabel metal2 s -150 5186 -150 5186 4 clk
port 6 nsew
rlabel metal2 s 8719 9296 8719 9296 4 men
port 7 nsew
flabel metal1 s 370 -345 370 -345 0 FreeSans 700 0 0 0 WEN
port 8 nsew
flabel metal3 s -311 -920 -311 -920 0 FreeSans 700 0 0 0 VSS
port 1 nsew
flabel metal3 s -311 -467 -311 -467 0 FreeSans 700 0 0 0 VDD
port 2 nsew
flabel metal3 s -311 132 -311 132 0 FreeSans 700 0 0 0 VDD
port 2 nsew
flabel metal3 s -311 1035 -311 1035 0 FreeSans 700 0 0 0 VSS
port 1 nsew
rlabel metal3 s 8856 3133 8856 3133 4 tblhl
port 3 nsew
flabel metal1 s 4631 812 4631 812 0 FreeSans 700 0 0 0 GWE
port 9 nsew
rlabel metal2 s 6127 -126 6127 -126 4 cen
port 5 nsew
<< properties >>
string path 25.525 19.160 25.525 21.230 
<< end >>
