magic
tech gf180mcuD
magscale 1 10
timestamp 1765480160
<< metal2 >>
rect -119 597 119 624
rect -119 -557 -93 597
rect 93 -557 119 597
rect -119 -584 119 -557
<< via2 >>
rect -93 -557 93 597
<< metal3 >>
rect -119 597 119 624
rect -119 -557 -93 597
rect 93 -557 119 597
rect -119 -584 119 -557
<< end >>
