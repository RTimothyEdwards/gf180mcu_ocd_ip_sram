magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< polysilicon >>
rect -41 211 14 245
rect 118 211 173 245
rect -41 -34 14 0
rect 118 -34 173 0
use nmos_5p04310591302039_256x8m81  nmos_5p04310591302039_256x8m81_0
timestamp 1763564386
transform 1 0 -14 0 1 0
box -116 -44 276 255
<< end >>
