magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal2 >>
rect -70 193 70 200
rect -70 -193 -63 193
rect 63 -193 70 193
rect -70 -200 70 -193
<< via2 >>
rect -63 -193 63 193
<< metal3 >>
rect -70 193 70 200
rect -70 -193 -63 193
rect 63 -193 70 193
rect -70 -200 70 -193
<< end >>
