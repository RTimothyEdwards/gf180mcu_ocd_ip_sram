magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nwell >>
rect -226 -219 1235 842
<< pmos >>
rect -46 236 455 749
rect 560 236 1061 749
<< pdiff >>
rect -140 735 -46 749
rect -140 249 -122 735
rect -76 249 -46 735
rect -140 236 -46 249
rect 455 735 560 749
rect 455 249 485 735
rect 531 249 560 735
rect 455 236 560 249
rect 1061 735 1149 749
rect 1061 249 1090 735
rect 1136 249 1149 735
rect 1061 236 1149 249
<< pdiffc >>
rect -122 249 -76 735
rect 485 249 531 735
rect 1090 249 1136 735
<< psubdiff >>
rect -126 988 1134 1001
rect -126 942 -62 988
rect 1071 942 1134 988
rect -126 928 1134 942
<< nsubdiff >>
rect -110 125 1118 138
rect -110 79 -62 125
rect 1071 79 1118 125
rect -110 36 1118 79
<< psubdiffcont >>
rect -62 942 1071 988
<< nsubdiffcont >>
rect -62 79 1071 125
<< polysilicon >>
rect -46 845 1061 858
rect -46 799 54 845
rect 1015 799 1061 845
rect -46 785 1061 799
rect -46 749 455 785
rect 560 749 1061 785
rect -46 191 455 236
rect 560 191 1061 236
<< polycontact >>
rect 54 799 1015 845
<< metal1 >>
rect -126 988 1134 1001
rect -126 942 -62 988
rect 1071 942 1134 988
rect -126 845 482 942
rect 534 845 1134 942
rect -126 799 54 845
rect 1015 799 1134 845
rect -126 795 1134 799
rect -130 735 -41 747
rect -130 619 -122 735
rect -76 619 -41 735
rect -130 271 -127 619
rect -71 271 -41 619
rect -130 249 -122 271
rect -76 249 -41 271
rect -130 238 -41 249
rect 450 735 567 748
rect 450 619 485 735
rect 531 619 567 735
rect 450 271 482 619
rect 534 271 567 619
rect 450 249 485 271
rect 531 249 567 271
rect 450 240 567 249
rect 451 236 567 240
rect 1055 735 1142 746
rect 1055 619 1090 735
rect 1136 619 1142 735
rect 1055 271 1085 619
rect 1141 271 1142 619
rect 1055 249 1090 271
rect 1136 249 1142 271
rect 1055 237 1142 249
rect -110 125 1118 138
rect -110 79 -62 125
rect 1071 79 1118 125
rect -110 36 1118 79
<< via1 >>
rect 482 942 534 973
rect 482 845 534 942
rect 482 822 534 845
rect -127 271 -122 619
rect -122 271 -76 619
rect -76 271 -71 619
rect 482 271 485 619
rect 485 271 531 619
rect 531 271 534 619
rect 1085 271 1090 619
rect 1090 271 1136 619
rect 1136 271 1141 619
<< metal2 >>
rect 471 973 545 987
rect 471 877 482 973
rect 534 877 545 973
rect 471 821 479 877
rect 537 821 545 877
rect 471 789 545 821
rect -135 621 1144 651
rect -135 269 -127 621
rect -71 619 1144 621
rect -71 271 482 619
rect 534 271 1085 619
rect 1141 271 1144 619
rect -71 269 1144 271
rect -135 240 1144 269
<< via2 >>
rect 479 822 482 877
rect 482 822 534 877
rect 534 822 537 877
rect 479 821 537 822
rect -127 619 -71 621
rect -127 271 -71 619
rect 1085 271 1141 619
rect -127 269 -71 271
<< metal3 >>
rect -150 621 -56 2597
rect -150 269 -127 621
rect -71 269 -56 621
rect -150 0 -56 269
rect 152 0 246 3737
rect 462 877 556 3808
rect 462 821 479 877
rect 537 821 556 877
rect 462 16 556 821
rect 770 16 864 3722
rect 1067 619 1161 2597
rect 1067 271 1085 619
rect 1141 271 1161 619
rect 1067 16 1161 271
<< end >>
