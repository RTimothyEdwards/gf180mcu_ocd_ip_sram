magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< nwell >>
rect -142 7186 550 8659
rect -4 6126 435 7186
rect -4 6086 436 6126
rect -3 5307 436 6086
rect -3 2035 436 2594
rect -3 1824 529 2035
rect -142 1381 529 1824
<< pmos >>
rect 96 7833 152 8152
rect 281 7833 337 8152
rect 96 7291 152 7610
rect 281 7291 337 7610
rect 64 1469 120 1608
rect 232 1469 288 1608
<< pdiff >>
rect -46 8139 96 8152
rect -46 7858 -23 8139
rect 23 7858 96 8139
rect -46 7833 96 7858
rect 152 8139 281 8152
rect 152 7858 193 8139
rect 240 7858 281 8139
rect 152 7833 281 7858
rect 337 8139 455 8152
rect 337 7858 367 8139
rect 413 7858 455 8139
rect 337 7833 455 7858
rect -46 7597 96 7610
rect -46 7316 -23 7597
rect 23 7316 96 7597
rect -46 7291 96 7316
rect 152 7597 281 7610
rect 152 7316 193 7597
rect 240 7316 281 7597
rect 152 7291 281 7316
rect 337 7597 455 7610
rect 337 7316 367 7597
rect 413 7316 455 7597
rect 337 7291 455 7316
rect -46 1577 64 1608
rect -46 1530 -23 1577
rect 23 1530 64 1577
rect -46 1469 64 1530
rect 120 1577 232 1608
rect 120 1530 154 1577
rect 200 1530 232 1577
rect 120 1469 232 1530
rect 288 1577 434 1608
rect 288 1530 329 1577
rect 375 1530 434 1577
rect 288 1469 434 1530
<< pdiffc >>
rect -23 7858 23 8139
rect 193 7858 240 8139
rect 367 7858 413 8139
rect -23 7316 23 7597
rect 193 7316 240 7597
rect 367 7316 413 7597
rect -23 1530 23 1577
rect 154 1530 200 1577
rect 329 1530 375 1577
<< nsubdiff >>
rect 0 8443 455 8555
rect 385 1885 434 1997
<< polysilicon >>
rect 96 8152 152 8362
rect 281 8152 337 8362
rect 96 7610 152 7833
rect 281 7610 337 7833
rect 96 7253 152 7291
rect 281 7253 337 7291
rect 96 7192 337 7253
rect 173 7009 229 7192
rect 175 5368 231 5469
rect 175 3767 231 4427
rect 175 3043 231 3194
rect 175 2982 244 2986
rect 175 2783 259 2847
rect 175 2726 231 2783
rect 64 1768 288 1837
rect 64 1608 120 1768
rect 232 1608 288 1768
rect 64 1295 120 1469
rect 232 1295 288 1469
<< metal1 >>
rect -40 8360 434 8558
rect -40 8139 102 8360
rect -40 7858 -23 8139
rect 23 7858 102 8139
rect -40 7597 102 7858
rect 176 8139 256 8304
rect 176 7858 193 8139
rect 240 7858 256 8139
rect 176 7840 256 7858
rect 330 8139 434 8360
rect 330 7858 367 8139
rect 413 7858 434 8139
rect -40 7316 -23 7597
rect 23 7316 102 7597
rect -40 7297 102 7316
rect 176 7597 256 7762
rect 176 7316 193 7597
rect 240 7316 256 7597
rect 176 7297 256 7316
rect 330 7597 434 7858
rect 330 7316 367 7597
rect 413 7316 434 7597
rect 330 7297 434 7316
rect 54 7189 317 7241
rect 40 6634 153 6760
rect 277 6634 390 6760
rect 49 5405 123 6027
rect 303 5405 384 6027
rect 49 5093 98 5405
rect 153 5355 280 5356
rect 153 5309 188 5355
rect 234 5345 280 5355
rect 153 5294 202 5309
rect 254 5294 280 5345
rect 153 5228 280 5294
rect 335 5093 384 5405
rect 49 4459 128 5093
rect 260 5080 384 5093
rect 306 4499 384 5080
rect 254 4389 384 4499
rect 31 4322 384 4389
rect -49 4020 434 4114
rect 33 3897 392 3965
rect 33 3097 131 3897
rect 33 2742 107 3097
rect 306 3091 384 3722
rect 168 2943 266 3038
rect 153 2792 280 2887
rect 328 2742 384 3091
rect 33 2096 126 2742
rect 304 2096 384 2742
rect -40 1899 40 1983
rect 371 1899 434 1983
rect -39 1577 39 1899
rect 95 1775 282 1843
rect 384 1671 434 1899
rect -39 1530 -23 1577
rect 23 1530 39 1577
rect -39 1499 39 1530
rect 136 1577 217 1671
rect 136 1530 154 1577
rect 200 1530 217 1577
rect -40 1164 39 1314
rect 136 1230 217 1530
rect 312 1577 434 1671
rect 312 1530 329 1577
rect 375 1530 434 1577
rect 312 1499 434 1530
rect 307 1164 434 1314
rect -40 1058 434 1164
<< metal2 >>
rect 53 8252 109 8659
rect 172 8360 261 8558
rect 53 8182 233 8252
rect 53 4459 109 8182
rect 344 7701 400 8659
rect 204 7632 400 7701
rect -107 1047 -46 4323
rect 209 3765 266 5356
rect 344 3878 400 7632
rect 56 3709 266 3765
rect 56 2873 112 3709
rect 175 2942 401 3010
rect 56 2865 176 2873
rect 56 2812 215 2865
rect 56 2805 176 2812
rect 56 1671 112 2805
rect 336 1843 401 2942
rect 266 1775 401 1843
rect 56 1614 186 1671
rect 172 1054 261 1205
<< metal3 >>
rect -45 7296 650 8615
rect 0 4064 651 5225
rect 0 3781 651 3931
rect 0 3536 650 3687
rect 0 3291 650 3441
rect 0 3056 650 3207
rect 0 2831 650 2981
rect 0 2581 650 2732
rect 0 2331 650 2481
rect 0 2091 650 2241
rect 0 1632 650 1941
rect 0 914 650 1232
use M1_NWELL$$46277676_512x8m81  M1_NWELL$$46277676_512x8m81_0
timestamp 1763765945
transform 1 0 217 0 1 8499
box -265 -159 265 159
use M1_NWELL$$47121452_512x8m81  M1_NWELL$$47121452_512x8m81_0
timestamp 1763765945
transform 1 0 165 0 1 1941
box -320 -159 320 159
use M1_PACTIVE4310591302075_512x8m81  M1_PACTIVE4310591302075_512x8m81_0
timestamp 1763765945
transform 1 0 170 0 1 1058
box -161 -36 161 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1763765945
transform 1 0 211 0 1 3012
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1763765945
transform 1 0 217 0 1 2818
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_2
timestamp 1763765945
transform 1 0 177 0 1 1808
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_3
timestamp 1763765945
transform 1 0 211 0 1 5332
box -36 -36 36 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_0
timestamp 1763765945
transform 1 0 212 0 1 7217
box -62 -36 62 36
use M1_PSUB$$45111340_512x8m81_0  M1_PSUB$$45111340_512x8m81_0_0
timestamp 1763765945
transform 1 0 0 0 1 4069
box -56 -58 56 58
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_0
timestamp 1763765945
transform 0 1 217 -1 0 2839
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_1
timestamp 1763765945
transform 1 0 67 0 1 6697
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_2
timestamp 1763765945
transform 1 0 230 0 1 7659
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_3
timestamp 1763765945
transform 1 0 203 0 1 8214
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_4
timestamp 1763765945
transform 1 0 73 0 1 5964
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_5
timestamp 1763765945
transform 1 0 178 0 1 1603
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_6
timestamp 1763765945
transform 1 0 228 0 1 5291
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_7
timestamp 1763765945
transform 1 0 364 0 1 6697
box -34 -63 34 63
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_0
timestamp 1763765945
transform 1 0 364 0 1 3934
box -35 -56 35 55
use M3_M2$$43368492_512x8m81_0  M3_M2$$43368492_512x8m81_0_0
timestamp 1763765945
transform 1 0 98 0 1 4143
box -45 -123 45 123
use nmos_5p0431059130200_512x8m81  nmos_5p0431059130200_512x8m81_0
timestamp 1763765945
transform 1 0 175 0 -1 5093
box -88 -44 144 679
use nmos_5p0431059130200_512x8m81  nmos_5p0431059130200_512x8m81_1
timestamp 1763765945
transform 1 0 175 0 -1 3726
box -88 -44 144 679
use nmos_5p0431059130202_512x8m81  nmos_5p0431059130202_512x8m81_0
timestamp 1763765945
transform 1 0 96 0 1 1232
box -124 -44 285 98
use pmos_5p0431059130201_512x8m81  pmos_5p0431059130201_512x8m81_0
timestamp 1763765945
transform 1 0 175 0 -1 2712
box -174 -86 230 721
use pmos_5p0431059130201_512x8m81  pmos_5p0431059130201_512x8m81_1
timestamp 1763765945
transform 1 0 173 0 -1 6977
box -174 -86 230 721
use pmos_5p0431059130201_512x8m81  pmos_5p0431059130201_512x8m81_2
timestamp 1763765945
transform 1 0 175 0 -1 6132
box -174 -86 230 721
use via1_2_512x8m81_0  via1_2_512x8m81_0_0
timestamp 1763765945
transform 1 0 184 0 1 1011
box 0 0 65 89
use via1_R90_512x8m81_0  via1_R90_512x8m81_0_0
timestamp 1763765945
transform 0 -1 264 1 0 2943
box 0 0 65 89
use via1_R90_512x8m81_0  via1_R90_512x8m81_0_1
timestamp 1763765945
transform 0 -1 261 1 0 8491
box 0 0 65 89
use via1_R90_512x8m81_0  via1_R90_512x8m81_0_2
timestamp 1763765945
transform 0 -1 261 1 0 8361
box 0 0 65 89
use via1_R270_512x8m81_0  via1_R270_512x8m81_0_0
timestamp 1763765945
transform 0 1 221 -1 0 1843
box 0 0 67 89
use via1_x2_R90_512x8m81_0  via1_x2_R90_512x8m81_0_0
timestamp 1763765945
transform 0 1 -107 1 0 4331
box -8 0 72 215
use via2_R90_512x8m81_0  via2_R90_512x8m81_0_0
timestamp 1763765945
transform 0 -1 261 1 0 8361
box 0 0 65 89
use via2_R90_512x8m81_0  via2_R90_512x8m81_0_1
timestamp 1763765945
transform 0 -1 261 1 0 8491
box 0 0 65 89
<< labels >>
rlabel metal2 s 362 8351 362 8351 4 b
port 3 nsew
rlabel metal2 s 73 8351 73 8351 4 bb
port 4 nsew
rlabel metal1 s 181 7190 181 7190 4 pcb
port 8 nsew
rlabel metal3 s 212 4328 212 4328 4 vss
port 1 nsew
rlabel metal3 s 222 8438 222 8438 4 vdd
port 2 nsew
rlabel metal1 s 222 1916 222 1916 4 vdd
port 2 nsew
rlabel metal2 s 199 1822 199 1822 4 ypass
port 6 nsew
rlabel metal1 s 344 1823 344 1823 4 d
port 7 nsew
rlabel metal2 s 0 1066 0 1066 4 db
port 5 nsew
rlabel metal3 s 189 1137 189 1137 4 vss
port 1 nsew
<< properties >>
string path 0.525 61.850 0.525 27.925 
<< end >>
