magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -44 713 44 731
rect -44 -713 -28 713
rect 28 -713 44 713
rect -44 -732 44 -713
<< via2 >>
rect -28 -713 28 713
<< metal3 >>
rect -45 713 45 732
rect -45 -713 -28 713
rect 28 -713 45 713
rect -45 -732 45 -713
<< end >>
