magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect 5024 6554 5936 7070
rect 4659 4844 8559 5394
rect 4713 2911 8559 4844
rect 4839 557 8346 1390
<< pmos >>
rect 5231 6653 5287 6865
rect 5367 6653 5423 6865
rect 5544 6653 5600 6865
rect 5673 6653 5729 6865
<< pdiff >>
rect 5119 6850 5231 6865
rect 5119 6678 5143 6850
rect 5189 6678 5231 6850
rect 5119 6653 5231 6678
rect 5287 6653 5367 6865
rect 5423 6850 5544 6865
rect 5423 6678 5457 6850
rect 5503 6678 5544 6850
rect 5423 6653 5544 6678
rect 5600 6653 5673 6865
rect 5729 6850 5840 6865
rect 5729 6678 5770 6850
rect 5817 6678 5840 6850
rect 5729 6653 5840 6678
<< pdiffc >>
rect 5143 6678 5189 6850
rect 5457 6678 5503 6850
rect 5770 6678 5817 6850
<< psubdiff >>
rect 5727 7588 8460 7622
rect 5727 7541 5793 7588
rect 8385 7541 8460 7588
rect 5727 7506 8460 7541
<< psubdiffcont >>
rect 5793 7541 8385 7588
<< polysilicon >>
rect 5203 7111 5259 7127
rect 5564 7126 5623 7332
rect 5231 6865 5287 7111
rect 5367 7081 5623 7126
rect 5367 7066 5600 7081
rect 5367 6865 5423 7066
rect 5544 6865 5600 7066
rect 5673 7014 5816 7072
rect 5673 7007 5751 7014
rect 5673 6865 5729 7007
rect 6327 6998 6383 7126
rect 6246 6944 6462 6998
rect 6246 6865 6302 6944
rect 6406 6865 6462 6944
rect 5231 6602 5287 6653
rect 5367 6602 5423 6653
rect 5544 6602 5600 6653
rect 5673 6602 5729 6653
<< metal1 >>
rect 4635 7588 8460 7616
rect 4635 7541 5793 7588
rect 8385 7541 8460 7588
rect 4635 7513 8460 7541
rect 5126 7173 5207 7513
rect 5282 7106 5364 7387
rect 5439 7173 5520 7513
rect 5282 7023 5520 7106
rect 5126 6850 5207 6943
rect 5126 6678 5143 6850
rect 5189 6678 5207 6850
rect 5126 6659 5207 6678
rect 5439 6850 5520 7023
rect 6241 7077 6323 7292
rect 6398 7221 6479 7511
rect 7115 7077 7205 7078
rect 6241 6984 7205 7077
rect 5439 6678 5457 6850
rect 5503 6678 5520 6850
rect 5439 6603 5520 6678
rect 5753 6895 5834 6943
rect 5753 6850 6240 6895
rect 5753 6678 5770 6850
rect 5817 6678 6240 6850
rect 6316 6731 6397 6984
rect 5753 6668 6240 6678
rect 6472 6668 6756 6895
rect 5753 6659 5834 6668
rect 5439 6519 6438 6603
rect 5393 3261 5474 3262
rect 5388 2879 5479 3261
<< metal2 >>
rect 503 7586 594 7679
rect 751 7586 841 7679
rect 1647 7586 1737 7679
rect 1900 7586 1991 7679
rect 2789 7586 2879 7679
rect 3036 7586 3127 7679
rect 3951 7586 4041 7679
rect 4177 7586 4267 7679
rect 5578 7357 5668 7451
rect 4984 7014 5846 7108
rect 5948 3982 6038 6603
rect 5588 3888 6038 3982
rect 5588 2853 5679 3888
rect 5748 2455 5838 3261
rect 6572 2738 6662 3261
rect 6932 2314 7022 3261
rect 7115 3187 7205 6974
rect 7756 2597 7846 3261
rect 8115 2173 8206 3099
rect 5786 148 5877 242
rect 6970 148 7060 242
rect 8154 148 8244 242
<< metal3 >>
rect 4753 7013 8515 7679
rect 0 6435 8515 6934
rect 0 5705 8550 6342
rect 0 3563 8563 5469
rect 0 1563 8389 2041
rect 0 754 8389 1390
rect 8225 366 8315 459
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_0
timestamp 1763476864
transform 1 0 3194 0 1 2772
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_1
timestamp 1763476864
transform 1 0 2723 0 1 2772
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_2
timestamp 1763476864
transform 1 0 280 0 1 2912
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_3
timestamp 1763476864
transform 1 0 1064 0 1 2912
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_4
timestamp 1763476864
transform 1 0 4024 0 1 2629
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_5
timestamp 1763476864
transform 1 0 4181 0 1 2205
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_6
timestamp 1763476864
transform 1 0 750 0 1 2205
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_7
timestamp 1763476864
transform 1 0 593 0 1 2629
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_8
timestamp 1763476864
transform 1 0 3350 0 1 2488
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_9
timestamp 1763476864
transform 1 0 2566 0 1 2488
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_10
timestamp 1763476864
transform 1 0 3867 0 1 2347
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_11
timestamp 1763476864
transform 1 0 4337 0 1 2347
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_12
timestamp 1763476864
transform 1 0 2050 0 1 2347
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_13
timestamp 1763476864
transform 1 0 1579 0 1 2347
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_14
timestamp 1763476864
transform 1 0 1893 0 1 2205
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_15
timestamp 1763476864
transform 1 0 1736 0 1 2629
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_16
timestamp 1763476864
transform 1 0 4494 0 1 2488
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_17
timestamp 1763476864
transform 1 0 2207 0 1 2912
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_18
timestamp 1763476864
transform 1 0 1423 0 1 2912
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_19
timestamp 1763476864
transform 1 0 3710 0 1 2488
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_20
timestamp 1763476864
transform 1 0 907 0 1 2772
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_21
timestamp 1763476864
transform 1 0 436 0 1 2772
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_22
timestamp 1763476864
transform 1 0 2880 0 1 2629
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_23
timestamp 1763476864
transform 1 0 3037 0 1 2205
box -67 -48 67 47
use M1_POLY2_R270_512x8m81  M1_POLY2_R270_512x8m81_0
timestamp 1763476864
transform 0 -1 5126 -1 0 7063
box -48 -123 48 123
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_0
timestamp 1763476864
transform 1 0 5600 0 1 7270
box -36 -126 60 122
use M1_POLY24310591302030_512x8m81  M1_POLY24310591302030_512x8m81_0
timestamp 1763476864
transform 1 0 6349 0 1 6583
box -95 -36 95 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1763476864
transform 1 0 5786 0 1 7043
box -36 -36 36 36
use M2_M1$$34864172_512x8m81  M2_M1$$34864172_512x8m81_0
timestamp 1763476864
transform -1 0 5103 0 1 7061
box -119 -46 119 46
use M2_M1$$34864172_512x8m81  M2_M1$$34864172_512x8m81_1
timestamp 1763476864
transform 1 0 5993 0 1 6556
box -119 -46 119 46
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1763476864
transform 1 0 5623 0 1 7328
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_1
timestamp 1763476864
transform 1 0 7160 0 1 6979
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_2
timestamp 1763476864
transform 1 0 5992 0 1 6804
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_3
timestamp 1763476864
transform 1 0 6711 0 1 6773
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_4
timestamp 1763476864
transform 1 0 5161 0 1 6763
box -43 -122 43 122
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_0
timestamp 1763476864
transform 1 0 6437 0 1 7363
box -44 -198 44 198
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_1
timestamp 1763476864
transform 1 0 5469 0 1 7403
box -44 -198 44 198
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_2
timestamp 1763476864
transform 1 0 5161 0 1 7403
box -44 -198 44 198
use M2_M1$$46894124_512x8m81  M2_M1$$46894124_512x8m81_0
timestamp 1763476864
transform -1 0 8161 0 1 2205
box -44 -46 45 46
use M2_M1$$46894124_512x8m81  M2_M1$$46894124_512x8m81_1
timestamp 1763476864
transform -1 0 7801 0 1 2629
box -44 -46 45 46
use M2_M1$$46894124_512x8m81  M2_M1$$46894124_512x8m81_2
timestamp 1763476864
transform -1 0 5793 0 1 2488
box -44 -46 45 46
use M2_M1$$46894124_512x8m81  M2_M1$$46894124_512x8m81_3
timestamp 1763476864
transform -1 0 6977 0 1 2347
box -44 -46 45 46
use M2_M1$$46894124_512x8m81  M2_M1$$46894124_512x8m81_4
timestamp 1763476864
transform -1 0 6617 0 1 2770
box -44 -46 45 46
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_0
timestamp 1763476864
transform 1 0 5747 0 1 7046
box -63 -34 63 34
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_0
timestamp 1763476864
transform 1 0 5992 0 1 6804
box -44 -123 44 123
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_1
timestamp 1763476864
transform 1 0 6711 0 1 6773
box -44 -123 44 123
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_2
timestamp 1763476864
transform 1 0 5161 0 1 6763
box -44 -123 44 123
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_0
timestamp 1763476864
transform 1 0 6437 0 1 7363
box -45 -198 45 198
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_1
timestamp 1763476864
transform 1 0 5469 0 1 7403
box -45 -198 45 198
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_2
timestamp 1763476864
transform 1 0 5161 0 1 7403
box -45 -198 45 198
use nmos_1p2$$47342636_512x8m81  nmos_1p2$$47342636_512x8m81_0
timestamp 1763476864
transform 1 0 6341 0 1 7165
box -102 -44 130 170
use nmos_5p04310591302056_512x8m81  nmos_5p04310591302056_512x8m81_0
timestamp 1763476864
transform 1 0 5363 0 1 7168
box -88 -44 144 222
use nmos_5p04310591302056_512x8m81  nmos_5p04310591302056_512x8m81_1
timestamp 1763476864
transform 1 0 5203 0 1 7168
box -88 -44 144 222
use pmos_1p2$$47109164_512x8m81  pmos_1p2$$47109164_512x8m81_0
timestamp 1763476864
transform 1 0 6288 0 1 6663
box -216 -86 348 245
use xpredec1_bot_512x8m81  xpredec1_bot_512x8m81_0
timestamp 1763476864
transform 1 0 7155 0 1 442
box -74 -442 1276 5964
use xpredec1_bot_512x8m81  xpredec1_bot_512x8m81_1
timestamp 1763476864
transform 1 0 4788 0 1 442
box -74 -442 1276 5964
use xpredec1_bot_512x8m81  xpredec1_bot_512x8m81_2
timestamp 1763476864
transform 1 0 5971 0 1 442
box -74 -442 1276 5964
use xpredec1_xa_512x8m81  xpredec1_xa_512x8m81_0
timestamp 1763476864
transform -1 0 3060 0 1 7450
box -100 -7451 774 228
use xpredec1_xa_512x8m81  xpredec1_xa_512x8m81_1
timestamp 1763476864
transform -1 0 4204 0 1 7450
box -100 -7451 774 228
use xpredec1_xa_512x8m81  xpredec1_xa_512x8m81_2
timestamp 1763476864
transform -1 0 1917 0 1 7450
box -100 -7451 774 228
use xpredec1_xa_512x8m81  xpredec1_xa_512x8m81_3
timestamp 1763476864
transform -1 0 773 0 1 7450
box -100 -7451 774 228
use xpredec1_xa_512x8m81  xpredec1_xa_512x8m81_4
timestamp 1763476864
transform 1 0 2874 0 1 7450
box -100 -7451 774 228
use xpredec1_xa_512x8m81  xpredec1_xa_512x8m81_5
timestamp 1763476864
transform 1 0 4018 0 1 7450
box -100 -7451 774 228
use xpredec1_xa_512x8m81  xpredec1_xa_512x8m81_6
timestamp 1763476864
transform 1 0 1731 0 1 7450
box -100 -7451 774 228
use xpredec1_xa_512x8m81  xpredec1_xa_512x8m81_7
timestamp 1763476864
transform 1 0 587 0 1 7450
box -100 -7451 774 228
<< labels >>
rlabel metal3 s 8399 6679 8399 6679 4 vdd
port 1 nsew
rlabel metal3 s 8399 5992 8399 5992 4 vss
port 2 nsew
rlabel metal3 s 8399 4515 8399 4515 4 vdd
port 1 nsew
rlabel metal3 s 8247 1117 8247 1117 4 vdd
port 1 nsew
rlabel metal3 s 8269 1802 8269 1802 4 vss
port 2 nsew
rlabel metal3 s 8269 412 8269 412 4 vss
port 2 nsew
rlabel metal3 s 8399 7389 8399 7389 4 vss
port 2 nsew
rlabel metal2 s 5832 195 5832 195 4 A[2]
port 3 nsew
rlabel metal2 s 5029 7065 5029 7065 4 men
port 4 nsew
rlabel metal2 s 548 7632 548 7632 4 x[7]
port 5 nsew
rlabel metal2 s 796 7632 796 7632 4 x[6]
port 6 nsew
rlabel metal2 s 1692 7632 1692 7632 4 x[5]
port 7 nsew
rlabel metal2 s 1946 7632 1946 7632 4 x[4]
port 8 nsew
rlabel metal2 s 2834 7632 2834 7632 4 x[3]
port 9 nsew
rlabel metal2 s 3082 7632 3082 7632 4 x[2]
port 10 nsew
rlabel metal2 s 3997 7632 3997 7632 4 x[1]
port 11 nsew
rlabel metal2 s 4222 7632 4222 7632 4 x[0]
port 12 nsew
rlabel metal2 s 7016 195 7016 195 4 A[1]
port 13 nsew
rlabel metal2 s 8199 195 8199 195 4 A[0]
port 14 nsew
rlabel metal2 s 5623 7401 5623 7401 4 clk
port 15 nsew
<< end >>
