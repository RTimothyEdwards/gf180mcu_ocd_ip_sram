magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect -210 -159 210 159
<< nsubdiff >>
rect -109 23 109 56
rect -109 -23 -78 23
rect 78 -23 109 23
rect -109 -56 109 -23
<< nsubdiffcont >>
rect -78 -23 78 23
<< metal1 >>
rect -95 23 95 42
rect -95 -23 -78 23
rect 78 -23 95 23
rect -95 -42 95 -23
<< end >>
