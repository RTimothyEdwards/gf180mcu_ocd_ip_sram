magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal2 >>
rect -200 627 200 634
rect -200 -627 -193 627
rect 193 -627 200 627
rect -200 -634 200 -627
<< via2 >>
rect -193 -627 193 627
<< metal3 >>
rect -200 627 200 634
rect -200 -627 -193 627
rect 193 -627 200 627
rect -200 -634 200 -627
<< end >>
