magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< metal2 >>
rect -330 106 330 113
rect -330 -106 -323 106
rect 323 -106 330 106
rect -330 -113 330 -106
<< via2 >>
rect -323 -106 323 106
<< metal3 >>
rect -330 106 330 113
rect -330 -106 -323 106
rect 323 -106 330 106
rect -330 -113 330 -106
<< end >>
