magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< psubdiff >>
rect -284 23 284 37
rect -284 -23 -252 23
rect 252 -23 284 23
rect -284 -36 284 -23
<< psubdiffcont >>
rect -252 -23 252 23
<< metal1 >>
rect -270 23 270 37
rect -270 -23 -252 23
rect 252 -23 270 23
rect -270 -35 270 -23
<< end >>
