magic
tech gf180mcuD
magscale 1 10
timestamp 1765833632
<< error_s >>
rect 605 8003 645 8005
rect 1885 8003 1925 8005
<< nwell >>
rect 2849 7137 3760 7148
rect 2644 7040 3760 7137
rect 2644 6683 4661 7040
rect 2644 6674 3760 6683
rect 2512 5770 2834 5865
rect 2512 5688 2972 5770
rect 2512 5247 2966 5688
rect 2512 5234 2999 5247
rect 2507 3907 2999 5234
rect 3728 5233 3878 5741
rect 3728 3963 3877 5233
rect 4176 3963 4923 5302
rect 3802 2179 3848 2797
<< pmos >>
rect 3035 6773 3091 6933
rect 3195 6773 3251 6933
rect 3360 6773 3416 6933
rect 3497 6773 3553 6933
<< pdiff >>
rect 2944 6919 3035 6933
rect 2944 6798 2958 6919
rect 3004 6798 3035 6919
rect 2944 6773 3035 6798
rect 3091 6773 3195 6933
rect 3251 6919 3360 6933
rect 3251 6798 3280 6919
rect 3326 6798 3360 6919
rect 3251 6773 3360 6798
rect 3416 6773 3497 6933
rect 3553 6919 3665 6933
rect 3553 6798 3595 6919
rect 3642 6798 3665 6919
rect 3553 6773 3665 6798
<< pdiffc >>
rect 2958 6798 3004 6919
rect 3280 6798 3326 6919
rect 3595 6798 3642 6919
<< polysilicon >>
rect 3420 7357 3479 7444
rect 3035 6933 3091 7259
rect 3195 7246 3251 7259
rect 3390 7246 3449 7327
rect 3195 7171 3449 7246
rect 3195 6933 3251 7171
rect 3360 7164 3449 7171
rect 3360 6933 3416 7164
rect 3556 7096 3692 7155
rect 3497 7054 3692 7096
rect 3497 6933 3553 7054
rect 4151 7038 4207 7263
rect 4073 6984 4289 7038
rect 4073 6932 4129 6984
rect 4233 6932 4289 6984
rect 3035 6722 3091 6773
rect 3195 6722 3251 6773
rect 3360 6722 3416 6773
rect 3497 6722 3553 6773
rect 4073 6670 4129 6747
rect 4233 6670 4289 6748
<< metal1 >>
rect 2950 7920 3032 7975
rect 2950 7288 3031 7920
rect 3107 7226 3188 7421
rect 3264 7288 3345 7979
rect 4223 7920 4305 8003
rect 4223 7682 4304 7920
rect 3107 7143 3345 7226
rect 4076 7204 4123 7374
rect 4223 7341 4305 7682
rect 2950 6919 3031 7015
rect 2950 6798 2958 6919
rect 3004 6798 3031 6919
rect 2950 6779 3031 6798
rect 3264 6919 3345 7143
rect 3562 7075 3675 7146
rect 4076 7110 5013 7204
rect 3264 6798 3280 6919
rect 3326 6798 3345 6919
rect 3264 6723 3345 6798
rect 3577 6919 4041 7015
rect 3577 6798 3595 6919
rect 3642 6798 4041 6919
rect 4157 6851 4204 7110
rect 3577 6783 4041 6798
rect 4322 6788 4581 7015
rect 3577 6779 3658 6783
rect 3264 6639 4279 6723
rect 2557 5572 2806 5655
rect 3211 3941 3302 4323
<< metal2 >>
rect 457 7739 548 7833
rect 706 7739 797 7833
rect 1710 7739 1801 7833
rect 1963 7739 2054 7833
rect 3402 7477 3493 7571
rect 2809 7134 3675 7228
rect 3773 6630 3864 6723
rect 3773 4931 3863 6630
rect 3413 4838 3863 4931
rect 3413 3792 3503 4838
rect 3573 3772 3663 4714
rect 4397 3634 4487 4299
rect 4757 3492 4847 4724
rect 4929 2981 5020 7101
rect 3612 1858 3702 1952
rect 4795 1858 4886 1952
<< metal3 >>
rect -202 7203 5166 7784
rect -202 6605 5166 7066
rect -202 5963 5166 6542
rect -202 4385 5166 5869
rect 289 2787 5166 3265
rect 289 2340 5166 2705
rect 289 1814 5166 2267
use M1_NACTIVE4310591302028_3v256x8m81  M1_NACTIVE4310591302028_3v256x8m81_0
timestamp 1765833244
transform 1 0 2793 0 1 6896
box -122 -181 122 181
use M1_NACTIVE4310591302028_3v256x8m81  M1_NACTIVE4310591302028_3v256x8m81_1
timestamp 1765833244
transform 1 0 4537 0 1 6896
box -122 -181 122 181
use M1_PACTIVE_02_3v256x8m81  M1_PACTIVE_02_3v256x8m81_0
timestamp 1763766357
transform 1 0 3836 0 1 7963
box -1382 -56 1408 56
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_0
timestamp 1765833244
transform 1 0 2324 0 1 3818
box -67 -48 67 47
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_1
timestamp 1765833244
transform 1 0 1065 0 1 3961
box -67 -48 67 47
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_2
timestamp 1765833244
transform 1 0 1443 0 1 3818
box -67 -48 67 47
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_3
timestamp 1765833244
transform 1 0 2163 0 1 3535
box -67 -48 67 47
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_4
timestamp 1765833244
transform 1 0 345 0 1 3675
box -67 -48 67 47
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_5
timestamp 1765833244
transform 1 0 868 0 1 3535
box -67 -48 67 47
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_6
timestamp 1765833244
transform 1 0 179 0 1 3961
box -67 -48 67 47
use M1_POLY2$$44753964_3v256x8m81  M1_POLY2$$44753964_3v256x8m81_7
timestamp 1765833244
transform 1 0 1605 0 1 3675
box -67 -48 67 47
use M1_POLY24310591302019_3v256x8m81  M1_POLY24310591302019_3v256x8m81_0
timestamp 1765833244
transform 0 -1 2969 1 0 7175
box -36 -80 36 78
use M1_POLY24310591302019_3v256x8m81  M1_POLY24310591302019_3v256x8m81_1
timestamp 1765833244
transform 0 -1 3619 1 0 7091
box -36 -80 36 78
use M1_POLY24310591302019_3v256x8m81  M1_POLY24310591302019_3v256x8m81_2
timestamp 1765833244
transform 1 0 3449 0 1 7382
box -36 -80 36 78
use M1_POLY24310591302030_3v256x8m81  M1_POLY24310591302030_3v256x8m81_0
timestamp 1765833244
transform 1 0 4189 0 1 6706
box -95 -36 95 36
use M2_M1$$34864172_3v256x8m81  M2_M1$$34864172_3v256x8m81_0
timestamp 1763766357
transform 1 0 3818 0 1 6676
box -119 -46 119 46
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_0
timestamp 1765833244
transform 1 0 4975 0 1 7105
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_1
timestamp 1765833244
transform 1 0 2986 0 1 6883
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_2
timestamp 1765833244
transform 1 0 4536 0 1 6893
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_3
timestamp 1765833244
transform 1 0 2793 0 1 6883
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_4
timestamp 1765833244
transform 1 0 3448 0 1 7448
box -43 -122 43 122
use M2_M1$$43375660_R90_3v256x8m81  M2_M1$$43375660_R90_3v256x8m81_0
timestamp 1765833244
transform 0 -1 3819 1 0 6842
box -46 -119 46 119
use M2_M1$$43380780_3v256x8m81  M2_M1$$43380780_3v256x8m81_0
timestamp 1763766357
transform 1 0 2986 0 1 7523
box -44 -198 44 198
use M2_M1$$43380780_3v256x8m81  M2_M1$$43380780_3v256x8m81_1
timestamp 1763766357
transform 1 0 3294 0 1 7523
box -44 -198 44 198
use M2_M1$$43380780_3v256x8m81  M2_M1$$43380780_3v256x8m81_2
timestamp 1763766357
transform 1 0 4263 0 1 7483
box -44 -198 44 198
use M2_M1$$46894124_3v256x8m81  M2_M1$$46894124_3v256x8m81_0
timestamp 1765833244
transform 1 0 3618 0 1 3818
box -44 -46 45 46
use M2_M1$$46894124_3v256x8m81  M2_M1$$46894124_3v256x8m81_1
timestamp 1765833244
transform 1 0 4442 0 1 3677
box -44 -46 45 46
use M2_M1$$46894124_3v256x8m81  M2_M1$$46894124_3v256x8m81_2
timestamp 1765833244
transform 1 0 4802 0 1 3535
box -44 -46 45 46
use M2_M1431059130200_3v256x8m81  M2_M1431059130200_3v256x8m81_0
timestamp 1765833244
transform 1 0 2963 0 1 7173
box -63 -34 63 34
use M2_M1431059130200_3v256x8m81  M2_M1431059130200_3v256x8m81_1
timestamp 1765833244
transform 1 0 3612 0 1 7173
box -63 -34 63 34
use M3_M2$$43368492_R90_3v256x8m81  M3_M2$$43368492_R90_3v256x8m81_0
timestamp 1765833244
transform 0 -1 3819 1 0 6842
box -46 -119 46 119
use M3_M2$$47108140_3v256x8m81  M3_M2$$47108140_3v256x8m81_0
timestamp 1763766357
transform 1 0 2986 0 1 6807
box -45 -198 45 198
use M3_M2$$47108140_3v256x8m81  M3_M2$$47108140_3v256x8m81_1
timestamp 1763766357
transform 1 0 4536 0 1 6816
box -45 -198 45 198
use M3_M2$$47108140_3v256x8m81  M3_M2$$47108140_3v256x8m81_2
timestamp 1763766357
transform 1 0 2986 0 1 7523
box -45 -198 45 198
use M3_M2$$47108140_3v256x8m81  M3_M2$$47108140_3v256x8m81_3
timestamp 1763766357
transform 1 0 3294 0 1 7523
box -45 -198 45 198
use M3_M2$$47108140_3v256x8m81  M3_M2$$47108140_3v256x8m81_4
timestamp 1763766357
transform 1 0 2793 0 1 6807
box -45 -198 45 198
use M3_M2$$47108140_3v256x8m81  M3_M2$$47108140_3v256x8m81_5
timestamp 1763766357
transform 1 0 4263 0 1 7483
box -45 -198 45 198
use nmos_1p2$$46563372_3v256x8m81  nmos_1p2$$46563372_3v256x8m81_0
timestamp 1765833452
transform 1 0 4165 0 1 7285
box -102 -44 130 133
use nmos_5p04310591302040_3v256x8m81  nmos_5p04310591302040_3v256x8m81_0
timestamp 1765833244
transform 1 0 3035 0 1 7288
box -88 -44 144 171
use nmos_5p04310591302040_3v256x8m81  nmos_5p04310591302040_3v256x8m81_1
timestamp 1765833244
transform 1 0 3195 0 1 7288
box -88 -44 144 171
use pmos_5p04310591302069_3v256x8m81  pmos_5p04310591302069_3v256x8m81_0
timestamp 1763766357
transform 1 0 4101 0 1 6783
box -202 -86 362 192
use xpredec0_bot_3v256x8m81  xpredec0_bot_3v256x8m81_0
timestamp 1765833452
transform 1 0 3796 0 1 569
box -74 1247 1270 5997
use xpredec0_bot_3v256x8m81  xpredec0_bot_3v256x8m81_1
timestamp 1765833452
transform 1 0 2613 0 1 569
box -74 1247 1270 5997
use xpredec0_xa_3v256x8m81  xpredec0_xa_3v256x8m81_0
timestamp 1765833632
transform -1 0 2817 0 1 23
box 107 1783 1129 7982
use xpredec0_xa_3v256x8m81  xpredec0_xa_3v256x8m81_1
timestamp 1765833632
transform -1 0 1537 0 1 23
box 107 1783 1129 7982
use xpredec0_xa_3v256x8m81  xpredec0_xa_3v256x8m81_2
timestamp 1765833632
transform 1 0 947 0 1 23
box 107 1783 1129 7982
use xpredec0_xa_3v256x8m81  xpredec0_xa_3v256x8m81_3
timestamp 1765833632
transform 1 0 -333 0 1 23
box 107 1783 1129 7982
<< labels >>
rlabel metal2 s 2006 7786 2006 7786 4 x[0]
port 5 nsew
rlabel metal2 s 1752 7786 1752 7786 4 x[1]
port 6 nsew
rlabel metal2 s 751 7786 751 7786 4 x[2]
port 7 nsew
rlabel metal2 s 502 7786 502 7786 4 x[3]
port 8 nsew
rlabel metal2 s 3448 7521 3448 7521 4 clk
port 10 nsew
rlabel metal2 s 2854 7185 2854 7185 4 men
port 4 nsew
rlabel metal3 s 5068 6945 5068 6945 4 vdd
port 1 nsew
rlabel metal3 s 5068 7628 5068 7628 4 vss
port 2 nsew
rlabel metal3 s 5068 6210 5068 6210 4 vss
port 2 nsew
rlabel metal3 s 5068 4895 5068 4895 4 vdd
port 1 nsew
rlabel metal2 s 3654 1905 3654 1905 4 A[1]
port 9 nsew
rlabel metal2 s 4837 1905 4837 1905 4 A[0]
port 3 nsew
rlabel metal3 s 10233 3009 10233 3009 4 vss
port 2 nsew
rlabel metal3 s 5068 3009 5068 3009 4 vss
port 2 nsew
rlabel metal3 s 10233 2376 10233 2376 4 vdd
port 1 nsew
rlabel metal3 s 5068 2376 5068 2376 4 vdd
port 1 nsew
rlabel metal3 s 10233 1922 10233 1922 4 vss
port 2 nsew
rlabel metal3 s 5068 1922 5068 1922 4 vss
port 2 nsew
<< end >>
