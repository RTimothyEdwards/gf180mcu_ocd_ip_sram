magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< nwell >>
rect 798 5267 1239 5500
rect -134 3584 -130 5026
rect 217 4720 1239 5267
rect 265 4380 1239 4720
rect 798 3621 1239 4380
rect 1032 3571 1239 3621
rect 1332 1623 1669 1635
rect 208 1505 1669 1623
rect 208 1479 1824 1505
rect -156 926 1824 1479
rect 207 925 806 926
rect 1383 925 1824 926
rect 208 868 806 925
rect 1384 698 1824 925
<< nmos >>
rect 522 5417 578 5524
<< pmos >>
rect 451 5030 507 5169
rect 614 5030 670 5169
<< ndiff >>
rect 406 5476 522 5524
rect 406 5430 437 5476
rect 483 5430 522 5476
rect 406 5417 522 5430
rect 578 5476 684 5524
rect 578 5430 621 5476
rect 667 5430 684 5476
rect 578 5417 684 5430
<< pdiff >>
rect 340 5095 451 5169
rect 340 5049 357 5095
rect 403 5049 451 5095
rect 340 5030 451 5049
rect 507 5095 614 5169
rect 507 5049 539 5095
rect 585 5049 614 5095
rect 507 5030 614 5049
rect 670 5095 781 5169
rect 670 5049 719 5095
rect 765 5049 781 5095
rect 670 5030 781 5049
<< ndiffc >>
rect 437 5430 483 5476
rect 621 5430 667 5476
<< pdiffc >>
rect 357 5049 403 5095
rect 539 5049 585 5095
rect 719 5049 765 5095
<< polysilicon >>
rect 522 5524 578 5575
rect 522 5316 578 5417
rect 451 5218 670 5316
rect 451 5169 507 5218
rect 614 5169 670 5218
rect 451 4980 507 5030
rect 614 4980 670 5030
rect 497 4708 633 4855
rect 357 4666 727 4708
rect 357 4344 413 4666
rect 671 4344 727 4666
rect 44 3372 100 3640
rect 997 3614 1053 3635
rect 908 3519 1053 3614
rect 997 3398 1053 3519
rect 357 2191 727 2255
rect 44 2035 100 2054
rect 966 2034 1050 2101
rect 976 2030 1032 2034
rect 976 1796 1032 1862
rect 976 1754 1193 1796
rect 471 1604 527 1743
rect 976 1698 1032 1754
rect 1136 1696 1192 1754
rect 401 1561 617 1604
rect 401 1291 457 1378
rect 767 1306 1197 1348
rect 387 1250 471 1291
rect 387 1208 1037 1250
rect 981 1152 1037 1208
rect 1141 1155 1197 1306
rect 1533 1258 1589 1800
rect 419 890 475 945
rect 194 848 475 890
rect 194 847 329 848
rect 419 793 475 848
rect 579 792 635 950
rect 981 927 1036 998
rect 981 884 1179 927
rect 795 794 1019 829
rect 795 787 963 794
rect 1123 790 1179 884
<< metal1 >>
rect 248 6117 1446 6185
rect 248 5971 1446 6038
rect 31 5796 1446 5892
rect 114 5647 1106 5714
rect 413 5536 825 5587
rect 413 5476 494 5536
rect -32 4761 16 5469
rect 413 5430 437 5476
rect 483 5430 494 5476
rect 413 5424 494 5430
rect 562 5476 678 5488
rect 562 5430 621 5476
rect 667 5430 678 5476
rect 562 5387 678 5430
rect 326 5222 507 5315
rect 562 5163 612 5387
rect 346 5095 414 5154
rect 346 5049 357 5095
rect 403 5049 414 5095
rect 346 5036 414 5049
rect 531 5095 612 5163
rect 531 5049 539 5095
rect 585 5049 612 5095
rect 531 5036 612 5049
rect 363 4725 414 5036
rect 562 4781 612 5036
rect 694 5095 775 5163
rect 694 5082 719 5095
rect 694 5049 718 5082
rect 765 5049 775 5095
rect 694 5036 775 5049
rect 694 4725 744 5036
rect 1081 4727 1128 5445
rect 363 4673 744 4725
rect 278 4276 335 4404
rect 588 4274 645 4402
rect 116 3608 197 3863
rect 429 3608 511 3863
rect 923 3760 973 3863
rect 743 3676 973 3760
rect 116 3524 877 3608
rect -31 3197 19 3250
rect 116 3208 197 3524
rect 274 3317 334 3374
rect 429 3285 511 3524
rect 923 3460 973 3676
rect 754 3404 973 3460
rect 591 3336 651 3378
rect 754 3306 814 3404
rect 923 3295 973 3404
rect 1396 3359 1508 5422
rect 1057 2337 1508 3359
rect 432 2179 634 2246
rect 251 2039 1512 2123
rect 251 2019 332 2039
rect 37 1935 332 2019
rect 577 1645 627 1862
rect 486 1593 836 1645
rect 486 1424 536 1593
rect 158 1209 443 1285
rect 135 827 286 911
rect 340 895 391 1020
rect 340 843 590 895
rect -7 612 53 718
rect 340 692 391 843
rect 490 612 540 690
rect -7 560 540 612
rect 684 612 734 1056
rect 785 854 836 1593
rect 889 1348 970 1618
rect 900 1347 966 1348
rect 1045 1292 1127 1953
rect 1202 1348 1283 1518
rect 1045 1208 1283 1292
rect 780 779 840 854
rect 888 612 934 1091
rect 684 560 934 612
rect 1081 613 1128 1076
rect 1202 662 1283 1208
rect 1458 1144 1512 2039
rect 1648 1900 1669 2030
rect 1648 1814 1725 1900
rect 1669 1684 1725 1814
rect 1618 1039 1707 1255
rect 1539 613 1590 719
rect 1081 562 1590 613
<< metal2 >>
rect 277 3150 343 6185
rect 558 6044 621 6304
rect 558 5961 658 6044
rect 436 2183 501 5892
rect 592 3145 658 5961
rect 803 5579 869 6415
rect 1052 6117 1115 6264
rect 1463 5971 1525 6301
rect 752 5511 869 5579
rect 752 5355 818 5511
rect 767 741 833 1869
rect 485 673 833 741
<< metal3 >>
rect -32 3630 1719 5535
rect -32 1573 1719 3430
rect -32 946 1719 1448
use M1_NWELL08_3v1024x8m81  M1_NWELL08_3v1024x8m81_0
timestamp 1764525316
transform 1 0 0 0 1 1262
box -154 -216 154 216
use M1_NWELL4310591302032_3v1024x8m81  M1_NWELL4310591302032_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1021 0 1 5408
box -126 -85 127 87
use M1_PACTIVE4310591302027_3v1024x8m81  M1_PACTIVE4310591302027_3v1024x8m81_0
timestamp 1764525316
transform 1 0 23 0 1 694
box -53 -62 53 62
use M1_POLY24310591302031_3v1024x8m81  M1_POLY24310591302031_3v1024x8m81_0
timestamp 1764525316
transform 1 0 473 0 1 2219
box -36 -36 36 36
use M1_POLY24310591302031_3v1024x8m81  M1_POLY24310591302031_3v1024x8m81_1
timestamp 1764525316
transform 1 0 810 0 1 816
box -36 -36 36 36
use M1_POLY24310591302031_3v1024x8m81  M1_POLY24310591302031_3v1024x8m81_2
timestamp 1764525316
transform 1 0 1559 0 1 706
box -36 -36 36 36
use M1_POLY24310591302031_3v1024x8m81  M1_POLY24310591302031_3v1024x8m81_3
timestamp 1764525316
transform 1 0 1008 0 1 2071
box -36 -36 36 36
use M1_PSUB$$45111340_3v1024x8m81  M1_PSUB$$45111340_3v1024x8m81_0
timestamp 1764525316
transform 1 0 0 0 1 1703
box -56 -58 56 58
use M1_PSUB$$46892076_3v1024x8m81  M1_PSUB$$46892076_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1446 0 1 4177
box -56 -1771 56 1241
use M1_PSUB$$46892076_3v1024x8m81  M1_PSUB$$46892076_3v1024x8m81_1
timestamp 1764525316
transform 1 0 1446 0 1 4177
box -56 -1771 56 1241
use M1_PSUB$$46893100_3v1024x8m81  M1_PSUB$$46893100_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1335 0 1 3149
box -56 -742 56 203
use M1_PSUB$$46893100_3v1024x8m81  M1_PSUB$$46893100_3v1024x8m81_1
timestamp 1764525316
transform 1 0 1335 0 1 3149
box -56 -742 56 203
use M2_M1$$43375660_R90_3v1024x8m81  M2_M1$$43375660_R90_3v1024x8m81_0
timestamp 1764525316
transform 0 -1 73 1 0 1700
box -46 -119 46 119
use M2_M1$$46894124_3v1024x8m81  M2_M1$$46894124_3v1024x8m81_0
timestamp 1764525316
transform 1 0 469 0 1 5846
box -44 -46 45 46
use M3_M2$$43368492_R90_3v1024x8m81  M3_M2$$43368492_R90_3v1024x8m81_0
timestamp 1764525316
transform 0 -1 73 1 0 1700
box -46 -119 46 119
use M3_M2$$46895148_3v1024x8m81  M3_M2$$46895148_3v1024x8m81_0
timestamp 1764525316
transform 1 0 469 0 1 5846
box -45 -46 45 46
use nmos_1p2$$46563372_3v1024x8m81  nmos_1p2$$46563372_3v1024x8m81_0
timestamp 1764525316
transform 1 0 990 0 -1 1989
box -102 -44 130 133
use nmos_1p2$$46563372_3v1024x8m81  nmos_1p2$$46563372_3v1024x8m81_1
timestamp 1764525316
transform 1 0 485 0 1 1784
box -102 -44 130 133
use nmos_1p2$$46883884_3v1024x8m81  nmos_1p2$$46883884_3v1024x8m81_0
timestamp 1764525316
transform 1 0 685 0 1 2297
box -102 -44 130 1102
use nmos_1p2$$46883884_3v1024x8m81  nmos_1p2$$46883884_3v1024x8m81_1
timestamp 1764525316
transform 1 0 1011 0 1 2297
box -102 -44 130 1102
use nmos_1p2$$46883884_3v1024x8m81  nmos_1p2$$46883884_3v1024x8m81_2
timestamp 1764525316
transform 1 0 371 0 1 2297
box -102 -44 130 1102
use nmos_1p2$$46884908_3v1024x8m81  nmos_1p2$$46884908_3v1024x8m81_0
timestamp 1764525316
transform 1 0 58 0 1 2090
box -102 -44 130 1314
use nmos_5p04310591302010_3v1024x8m81  nmos_5p04310591302010_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1533 0 -1 2049
box -88 -44 144 255
use nmos_5p04310591302011_3v1024x8m81  nmos_5p04310591302011_3v1024x8m81_0
timestamp 1764525316
transform 1 0 447 0 -1 770
box -116 -44 276 133
use nmos_5p04310591302011_3v1024x8m81  nmos_5p04310591302011_3v1024x8m81_1
timestamp 1764525316
transform 1 0 991 0 1 661
box -116 -44 276 133
use pmos_1p2$$46273580_3v1024x8m81  pmos_1p2$$46273580_3v1024x8m81_0
timestamp 1764525316
transform 1 0 443 0 -1 1524
box -216 -86 348 192
use pmos_1p2$$46273580_3v1024x8m81  pmos_1p2$$46273580_3v1024x8m81_1
timestamp 1764525316
transform 1 0 1018 0 -1 1659
box -216 -86 348 192
use pmos_1p2$$46885932_3v1024x8m81  pmos_1p2$$46885932_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1023 0 1 1024
box -216 -86 348 175
use pmos_1p2$$46887980_3v1024x8m81  pmos_1p2$$46887980_3v1024x8m81_0
timestamp 1764525316
transform 1 0 58 0 1 3670
box -188 -86 216 1356
use pmos_1p2$$46889004_3v1024x8m81  pmos_1p2$$46889004_3v1024x8m81_0
timestamp 1764525316
transform 1 0 371 0 1 3670
box -188 -86 216 721
use pmos_1p2$$46889004_3v1024x8m81  pmos_1p2$$46889004_3v1024x8m81_1
timestamp 1764525316
transform 1 0 685 0 1 3670
box -188 -86 216 721
use pmos_5p0431059130201_3v1024x8m81  pmos_5p0431059130201_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1533 0 1 783
box -174 -86 230 721
use pmos_5p0431059130206_3v1024x8m81  pmos_5p0431059130206_3v1024x8m81_0
timestamp 1764525316
transform 1 0 447 0 1 967
box -202 -86 362 175
use pmos_5p0431059130209_3v1024x8m81  pmos_5p0431059130209_3v1024x8m81_0
timestamp 1764525316
transform 1 0 997 0 1 3670
box -174 -86 230 1144
use po_m1_3v1024x8m81  po_m1_3v1024x8m81_0
timestamp 1764525316
transform -1 0 638 0 -1 916
box -21 0 113 95
use po_m1_3v1024x8m81  po_m1_3v1024x8m81_1
timestamp 1764525316
transform 1 0 519 0 -1 4854
box -21 0 113 95
use po_m1_3v1024x8m81  po_m1_3v1024x8m81_2
timestamp 1764525316
transform 1 0 356 0 1 1208
box -21 0 113 95
use po_m1_3v1024x8m81  po_m1_3v1024x8m81_3
timestamp 1764525316
transform 1 0 32 0 1 1943
box -21 0 113 95
use po_m1_R90_3v1024x8m81  po_m1_R90_3v1024x8m81_0
timestamp 1764525316
transform 0 -1 897 1 0 3519
box 0 -21 95 113
use po_m1_R90_3v1024x8m81  po_m1_R90_3v1024x8m81_1
timestamp 1764525316
transform 0 -1 847 1 0 1306
box 0 -21 95 113
use po_m1_R270_3v1024x8m81  po_m1_R270_3v1024x8m81_0
timestamp 1764525316
transform 0 1 214 -1 0 916
box 0 -21 95 114
use po_m1_R270_3v1024x8m81  po_m1_R270_3v1024x8m81_1
timestamp 1764525316
transform 0 1 436 -1 0 5320
box 0 -21 95 114
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_0
timestamp 1764525316
transform -1 0 565 0 -1 1196
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_1
timestamp 1764525316
transform -1 0 702 0 -1 1440
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_2
timestamp 1764525316
transform -1 0 965 0 -1 1440
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_3
timestamp 1764525316
transform 1 0 -32 0 1 2686
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_4
timestamp 1764525316
transform 1 0 1057 0 1 2344
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_5
timestamp 1764525316
transform 1 0 -22 0 1 3029
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_6
timestamp 1764525316
transform 1 0 1057 0 1 3129
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_7
timestamp 1764525316
transform 1 0 1057 0 1 2686
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_8
timestamp 1764525316
transform 1 0 -32 0 1 1148
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_9
timestamp 1764525316
transform 1 0 402 0 1 1748
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_10
timestamp 1764525316
transform 1 0 1714 0 1 1040
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_11
timestamp 1764525316
transform 1 0 1066 0 1 3826
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_12
timestamp 1764525316
transform 1 0 -32 0 1 3826
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_13
timestamp 1764525316
transform 1 0 1066 0 1 4869
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_14
timestamp 1764525316
transform 1 0 -32 0 1 5265
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_15
timestamp 1764525316
transform 1 0 -32 0 1 4846
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_16
timestamp 1764525316
transform 1 0 1714 0 1 1685
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_17
timestamp 1764525316
transform 1 0 905 0 1 1748
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_18
timestamp 1764525316
transform 1 0 -32 0 1 2344
box -9 0 73 215
use via1_2_x2_3v1024x8m81  via1_2_x2_3v1024x8m81_19
timestamp 1764525316
transform 1 0 723 0 1 4939
box -9 0 73 215
use via1_2_x2_R90_3v1024x8m81  via1_2_x2_R90_3v1024x8m81_0
timestamp 1764525316
transform 0 -1 390 1 0 1374
box -9 0 73 215
use via1_2_x2_R90_3v1024x8m81  via1_2_x2_R90_3v1024x8m81_1
timestamp 1764525316
transform 0 -1 1128 1 0 5376
box -9 0 73 215
use via1_3v1024x8m81  via1_3v1024x8m81_0
timestamp 1764525316
transform 1 0 485 0 1 659
box 0 0 65 92
use via1_3v1024x8m81  via1_3v1024x8m81_1
timestamp 1764525316
transform 1 0 436 0 1 5222
box 0 0 65 92
use via1_R90_3v1024x8m81  via1_R90_3v1024x8m81_0
timestamp 1764525316
transform 0 -1 522 1 0 2179
box 0 0 65 89
use via1_x2_3v1024x8m81  via1_x2_3v1024x8m81_0
timestamp 1764525316
transform -1 0 1268 0 -1 1570
box -8 0 72 222
use via1_x2_3v1024x8m81  via1_x2_3v1024x8m81_1
timestamp 1764525316
transform 1 0 595 0 1 4387
box -8 0 72 222
use via1_x2_3v1024x8m81  via1_x2_3v1024x8m81_2
timestamp 1764525316
transform 1 0 277 0 1 4387
box -8 0 72 222
use via1_x2_3v1024x8m81  via1_x2_3v1024x8m81_3
timestamp 1764525316
transform 1 0 753 0 1 5355
box -8 0 72 222
use via1_x2_3v1024x8m81  via1_x2_3v1024x8m81_4
timestamp 1764525316
transform 1 0 280 0 1 3133
box -8 0 72 222
use via1_x2_3v1024x8m81  via1_x2_3v1024x8m81_5
timestamp 1764525316
transform 1 0 595 0 1 3133
box -8 0 72 222
use via1_x2_R90_3v1024x8m81  via1_x2_R90_3v1024x8m81_0
timestamp 1764525316
transform 0 -1 1610 1 0 5971
box -8 0 72 215
use via1_x2_R90_3v1024x8m81  via1_x2_R90_3v1024x8m81_1
timestamp 1764525316
transform 0 -1 1190 1 0 6117
box -8 0 72 215
use via1_x2_R90_3v1024x8m81  via1_x2_R90_3v1024x8m81_2
timestamp 1764525316
transform 0 -1 744 1 0 5971
box -8 0 72 215
use via1_x2_R90_3v1024x8m81  via1_x2_R90_3v1024x8m81_3
timestamp 1764525316
transform 0 -1 448 1 0 6117
box -8 0 72 215
use via2_x2_3v1024x8m81  via2_x2_3v1024x8m81_0
timestamp 1764525316
transform -1 0 1268 0 -1 1440
box -9 0 74 222
use via2_x2_3v1024x8m81  via2_x2_3v1024x8m81_1
timestamp 1764525316
transform 1 0 768 0 1 1647
box -9 0 74 222
<< labels >>
rlabel metal3 s 1040 4168 1040 4168 4 vdd
port 2 nsew
rlabel metal2 s 304 5597 304 5597 4 d
port 3 nsew
rlabel metal1 s 735 5854 735 5854 4 wep
port 6 nsew
rlabel metal1 s 877 6158 877 6158 4 d
port 3 nsew
rlabel metal1 s 975 6015 975 6015 4 db
port 4 nsew
rlabel metal2 s 829 5737 829 5737 4 vss
port 1 nsew
rlabel metal2 s 618 5597 618 5597 4 db
port 4 nsew
rlabel metal3 s 1089 2776 1089 2776 4 vss
port 1 nsew
rlabel metal1 s 263 875 263 875 4 datain
port 5 nsew
rlabel metal1 s 399 1259 399 1259 4 men
port 7 nsew
<< end >>
