magic
tech gf180mcuD
magscale 1 10
timestamp 1764700137
<< error_p >>
rect -75 0 -29 89
rect 85 0 131 89
<< nmos >>
rect 0 0 56 89
<< ndiff >>
rect -88 76 0 89
rect -88 13 -75 76
rect -29 13 0 76
rect -88 0 0 13
rect 56 76 144 89
rect 56 13 85 76
rect 131 13 144 76
rect 56 0 144 13
<< ndiffc >>
rect -75 13 -29 76
rect 85 13 131 76
<< polysilicon >>
rect 0 89 56 133
rect 0 -44 56 0
<< metal1 >>
rect -75 76 -29 89
rect -75 0 -29 13
rect 85 76 131 89
rect 85 0 131 13
<< labels >>
flabel ndiffc -40 44 -40 44 0 FreeSans 93 0 0 0 S
flabel ndiffc 96 44 96 44 0 FreeSans 93 0 0 0 D
<< end >>
