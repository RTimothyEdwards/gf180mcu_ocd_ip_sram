magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal2 >>
rect -1373 104 1373 123
rect -1373 -104 -1357 104
rect 1357 -104 1373 104
rect -1373 -122 1373 -104
<< via2 >>
rect -1357 -104 1357 104
<< metal3 >>
rect -1373 104 1373 123
rect -1373 -104 -1357 104
rect 1357 -104 1373 104
rect -1373 -123 1373 -104
<< end >>
