magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -330 1625 330 1632
rect -330 -1275 -323 1625
rect 323 -1275 330 1625
rect -330 -1282 330 -1275
<< via2 >>
rect -323 -1275 323 1625
<< metal3 >>
rect -330 1625 330 1632
rect -330 -1275 -323 1625
rect 323 -1275 330 1625
rect -330 -1282 330 -1275
<< end >>
