magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< metal1 >>
rect 2654 20538 4331 20632
rect 2837 17681 4185 17682
rect 2632 17546 4185 17681
<< metal2 >>
rect 2831 25266 3510 36851
rect 2831 4045 3531 25266
<< metal3 >>
rect 2338 25911 4138 26051
rect 2338 25784 3047 25911
rect 2338 25448 4138 25784
rect 2338 23755 4138 25160
rect 2338 22413 3531 23755
rect 2338 22214 4642 22413
rect 2338 20557 4445 21944
rect 2338 18459 3531 18849
rect 2338 18149 4445 18459
rect 2338 17432 4445 17750
rect 2338 17051 3047 17432
rect 2982 17050 3047 17051
rect 2338 14821 4445 16727
rect 2338 12769 4445 14621
rect 2338 12141 4445 12642
rect 2338 11770 3531 12141
rect 2338 11203 4445 11770
rect 2338 11183 3531 11203
rect 2338 9902 4445 10824
rect 2338 8484 4445 9438
rect 2338 7908 4445 8272
rect 2338 7842 3049 7908
rect 2338 7444 3047 7842
rect 2338 7141 4445 7444
rect 2338 6729 4445 7048
rect 2338 6338 3535 6729
rect 2338 6020 4445 6338
rect 2338 5572 4445 5818
rect 2338 5176 3037 5572
rect 2338 4929 4445 5176
rect 2338 4041 4445 4741
use M2_M14310591302080_3v1024x8m81  M2_M14310591302080_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2648 0 1 5374
box -113 -417 113 417
use M2_M14310591302080_3v1024x8m81  M2_M14310591302080_3v1024x8m81_1
timestamp 1764525316
transform 1 0 2648 0 1 10354
box -113 -417 113 417
use M2_M14310591302081_3v1024x8m81  M2_M14310591302081_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2648 0 1 17401
box -113 -330 113 330
use M2_M14310591302087_3v1024x8m81  M2_M14310591302087_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2648 0 1 25721
box -113 -243 113 243
use M2_M14310591302092_3v1024x8m81  M2_M14310591302092_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2648 0 1 13453
box -113 -655 113 1155
use M2_M14310591302093_3v1024x8m81  M2_M14310591302093_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2648 0 1 7789
box -113 -634 113 634
use M2_M14310591302093_3v1024x8m81  M2_M14310591302093_3v1024x8m81_1
timestamp 1764525316
transform 1 0 2648 0 1 20504
box -113 -634 113 634
use M3_M24310591302042_3v1024x8m81  M3_M24310591302042_3v1024x8m81_0
timestamp 1764525316
transform 1 0 3189 0 1 4388
box -330 -330 330 330
use M3_M24310591302042_3v1024x8m81  M3_M24310591302042_3v1024x8m81_1
timestamp 1764525316
transform 1 0 3189 0 1 18500
box -330 -330 330 330
use M3_M24310591302082_3v1024x8m81  M3_M24310591302082_3v1024x8m81_0
timestamp 1764525316
transform 1 0 3189 0 1 6579
box -330 -547 330 447
use M3_M24310591302083_3v1024x8m81  M3_M24310591302083_3v1024x8m81_0
timestamp 1764525316
transform 1 0 3189 0 1 23524
box -330 -1282 330 1632
use M3_M24310591302084_3v1024x8m81  M3_M24310591302084_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2648 0 1 13453
box -113 -655 113 1155
use M3_M24310591302085_3v1024x8m81  M3_M24310591302085_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2648 0 1 17401
box -113 -330 113 330
use M3_M24310591302086_3v1024x8m81  M3_M24310591302086_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2648 0 1 7789
box -113 -634 113 474
use M3_M24310591302086_3v1024x8m81  M3_M24310591302086_3v1024x8m81_1
timestamp 1764525316
transform 1 0 2648 0 1 21244
box -113 -634 113 474
use M3_M24310591302088_3v1024x8m81  M3_M24310591302088_3v1024x8m81_0
timestamp 1764525316
transform 1 0 3189 0 1 11910
box -330 -721 330 721
use M3_M24310591302089_3v1024x8m81  M3_M24310591302089_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2648 0 1 5374
box -113 -417 113 417
use M3_M24310591302089_3v1024x8m81  M3_M24310591302089_3v1024x8m81_1
timestamp 1764525316
transform 1 0 2648 0 1 10354
box -113 -417 113 417
use M3_M24310591302090_3v1024x8m81  M3_M24310591302090_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2648 0 1 25721
box -113 -243 113 243
use M3_M24310591302091_3v1024x8m81  M3_M24310591302091_3v1024x8m81_0
timestamp 1764525316
transform 1 0 3189 0 1 8965
box -330 -460 330 460
use M3_M24310591302094_3v1024x8m81  M3_M24310591302094_3v1024x8m81_0
timestamp 1764525316
transform 1 0 3189 0 1 15774
box -330 -938 330 938
<< end >>
