magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -118 257 119 275
rect -118 -257 -102 257
rect 102 -257 119 257
rect -118 -275 119 -257
<< via2 >>
rect -102 -257 102 257
<< metal3 >>
rect -119 257 119 275
rect -119 -257 -102 257
rect 102 -257 119 257
rect -119 -275 119 -257
<< end >>
