magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -44 1551 45 1570
rect -44 -1551 -28 1551
rect 28 -1551 45 1551
rect -44 -1570 45 -1551
<< via2 >>
rect -28 -1551 28 1551
<< metal3 >>
rect -45 1551 45 1570
rect -45 -1551 -28 1551
rect 28 -1551 45 1551
rect -45 -1570 45 -1551
<< end >>
