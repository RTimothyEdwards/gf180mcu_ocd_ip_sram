magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect -371 3355 531 3507
rect -371 2774 3558 3355
rect -371 1884 3622 2774
rect -371 436 -57 499
rect 2474 436 2915 437
rect 3393 436 3622 475
rect -371 38 3622 436
rect -371 -16 -44 38
<< polysilicon >>
rect 1589 3864 2442 3906
rect 116 3288 172 3616
rect 276 3288 332 3616
rect 753 3453 809 3475
rect 913 3453 969 3475
rect 1075 3453 1131 3475
rect 1235 3453 1291 3475
rect 1397 3453 1453 3460
rect 462 3411 1453 3453
rect 753 3190 809 3411
rect 913 3190 969 3411
rect 1074 3190 1130 3411
rect 1589 3340 1629 3864
rect 1742 3753 1798 3864
rect 1902 3753 1958 3864
rect 2064 3753 2120 3864
rect 2224 3753 2280 3864
rect 2386 3753 2442 3864
rect 2735 3383 2791 3468
rect 1234 3298 1629 3340
rect 1234 3190 1290 3298
rect 1409 3278 1629 3298
rect 1783 3331 2791 3383
rect 2895 3331 2951 3468
rect 3055 3331 3111 3468
rect 3215 3331 3271 3468
rect 1783 3288 3283 3331
rect 1409 3095 1572 3278
rect 1783 3155 1839 3288
rect 1943 3155 1999 3288
rect 2104 3155 2160 3288
rect 2264 3155 2320 3288
rect 2425 3155 2481 3288
rect 2585 3155 2641 3288
rect 2746 3155 2802 3288
rect 2906 3155 2962 3288
rect 3067 3155 3123 3288
rect 3227 3155 3283 3288
rect 116 2882 172 2893
rect 276 2882 332 2893
rect 116 2786 332 2882
rect 89 1924 145 2126
rect 249 1924 305 2126
rect 410 1924 466 2126
rect 570 1924 626 2126
rect 731 1924 787 2126
rect 891 1924 947 2126
rect 1052 1924 1108 2126
rect 1212 1924 1268 2126
rect 1373 1924 1429 2126
rect 1533 1924 1589 2126
rect 89 1881 1611 1924
rect 266 1650 322 1881
rect 428 1650 484 1881
rect 588 1650 644 1881
rect 750 1650 806 1881
rect 910 1650 966 1881
rect 1072 1650 1128 1881
rect 1232 1837 1611 1881
rect 1232 1650 1288 1837
rect 2010 1756 2066 2095
rect 1850 1700 2066 1756
rect 1850 1650 1906 1700
rect 2010 1648 2066 1700
rect 2171 1648 2227 2095
rect 2331 1648 2387 2095
rect 2636 1855 2692 2097
rect 2501 1853 2692 1855
rect 2797 1870 2853 2097
rect 2957 1870 3013 2095
rect 2797 1853 3013 1870
rect 2501 1827 3013 1853
rect 2501 1797 2856 1827
rect 2640 1647 2696 1797
rect 2800 1647 2856 1797
rect 1689 1103 1745 1310
rect 2171 1103 2227 1309
rect 1689 1061 2227 1103
rect 122 880 810 881
rect 115 879 810 880
rect 115 838 813 879
rect 115 747 171 838
rect 275 747 331 838
rect 436 747 492 838
rect 596 747 652 838
rect 757 747 813 838
rect 115 530 171 579
rect 275 530 331 579
rect 436 530 492 579
rect 596 530 652 579
rect 757 530 813 579
rect 115 433 186 530
rect 275 433 346 530
rect 436 433 507 530
rect 596 433 667 530
rect 757 433 828 530
rect 1149 529 1209 584
rect 940 470 1209 529
rect 130 336 186 433
rect 290 336 346 433
rect 451 336 507 433
rect 611 336 667 433
rect 772 336 828 433
rect 1153 355 1209 470
rect 1313 355 1369 578
rect 1656 570 1716 577
rect 1447 511 1716 570
rect 1660 359 1716 511
rect 1820 359 1876 577
rect 2153 527 2209 579
rect 1957 469 2213 527
rect 2321 495 2377 579
rect 2653 527 2709 578
rect 2157 358 2213 469
rect 2317 358 2373 495
rect 2446 469 2709 527
rect 2985 499 3041 533
rect 2653 383 2709 469
rect 2931 440 2975 499
rect 2985 440 3202 499
rect 2985 338 3041 440
rect 3145 336 3201 440
<< metal1 >>
rect 833 3871 2517 3917
rect 833 3815 913 3871
rect 201 3584 248 3749
rect 832 3687 913 3815
rect 1144 3601 1225 3871
rect 1458 3601 1539 3871
rect 1827 3601 1873 3871
rect 2149 3597 2195 3871
rect 2471 3659 2517 3871
rect 2804 3857 3198 3906
rect 201 3531 534 3584
rect 201 3236 248 3531
rect 483 3363 534 3531
rect 1667 3390 1713 3574
rect 1988 3390 2034 3572
rect 2310 3390 2356 3587
rect 830 3306 2356 3390
rect 830 3136 912 3306
rect 1144 3127 1225 3306
rect 2288 3294 2356 3306
rect 2288 3293 2345 3294
rect 1865 2812 1946 3050
rect 2177 2812 2258 3065
rect 2491 2812 2572 3065
rect 2804 2812 2886 3857
rect 3117 2812 3198 3857
rect 184 2747 729 2800
rect 1865 2744 3198 2812
rect 37 2604 1688 2688
rect 37 2327 119 2604
rect 323 2355 404 2604
rect 637 2355 717 2604
rect 981 2355 1062 2604
rect 1283 2355 1364 2604
rect 1607 2430 1688 2604
rect 166 1843 247 2251
rect 490 1843 570 2232
rect 813 1843 894 2220
rect 1136 1903 1218 2213
rect 1450 1903 1531 2335
rect 1136 1843 1531 1903
rect 166 1819 1531 1843
rect 166 1759 1218 1819
rect 1605 1808 1814 1918
rect 2077 1871 2158 2211
rect 2415 1871 2474 2196
rect 166 1530 247 1759
rect 490 1530 570 1759
rect 813 1530 894 1759
rect 1136 1530 1218 1759
rect 1920 1788 2558 1871
rect 353 1233 434 1530
rect 667 1233 747 1530
rect 980 1233 1061 1530
rect 1309 1233 1359 1424
rect 1920 1346 2002 1788
rect 2704 1513 2786 2206
rect 3024 1862 3100 2217
rect 353 1181 1359 1233
rect 604 1057 3129 1125
rect 3201 973 3468 1278
rect -261 877 3517 973
rect 851 740 1122 808
rect 211 533 260 680
rect 536 533 585 680
rect 851 533 900 740
rect 1070 577 1124 667
rect 1293 621 1341 812
rect 211 450 989 533
rect 211 231 260 450
rect 512 449 585 450
rect 826 449 900 450
rect 536 223 585 449
rect 854 233 900 449
rect 1078 248 1124 577
rect 1287 571 1347 621
rect 1400 618 1476 702
rect 1293 521 1341 571
rect 1425 248 1476 618
rect 1559 522 1610 684
rect 1559 474 1848 522
rect 1559 248 1610 474
rect 1933 248 1983 684
rect 2065 522 2116 684
rect 2406 600 2499 684
rect 2065 474 2355 522
rect 2065 242 2116 474
rect 2452 375 2499 600
rect 2421 242 2499 375
rect 2578 234 2625 673
rect 2593 233 2625 234
rect 3070 137 3120 685
<< metal2 >>
rect 602 1057 667 2816
rect 1437 2663 1502 3231
rect 1592 2797 1654 3383
rect 1592 2733 2006 2797
rect 1437 2595 1879 2663
rect 1943 2604 2006 2733
rect 1813 1730 1879 2595
rect 1144 1662 2296 1730
rect 1144 746 1210 1662
rect 3063 543 3129 1125
rect 3201 879 3468 1278
rect 1052 434 2792 501
<< metal3 >>
rect -250 3588 3587 3958
rect -252 2173 3500 3126
rect 2712 1918 2779 1919
rect 3028 1918 3093 1919
rect 1532 1851 3093 1918
rect -252 1353 3500 1782
rect -261 879 3517 1278
rect -252 502 3500 805
rect -252 88 3514 406
use M1_NWELL02_512x8m81  M1_NWELL02_512x8m81_0
timestamp 1763476864
transform 1 0 -217 0 -1 255
box -154 -159 154 159
use M1_NWELL03_512x8m81  M1_NWELL03_512x8m81_0
timestamp 1763476864
transform 1 0 3413 0 1 2329
box -210 -445 210 445
use M1_NWELL04_512x8m81  M1_NWELL04_512x8m81_0
timestamp 1763476864
transform 1 0 -217 0 1 2329
box -154 -445 154 445
use M1_PACTIVE4310591302034_512x8m81  M1_PACTIVE4310591302034_512x8m81_0
timestamp 1763476864
transform 1 0 -217 0 1 3762
box -36 -128 36 128
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_0
timestamp 1763476864
transform 1 0 688 0 1 919
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_1
timestamp 1763476864
transform 1 0 240 0 1 919
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_2
timestamp 1763476864
transform 1 0 224 0 1 2834
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_3
timestamp 1763476864
transform 1 0 530 0 1 3405
box -67 -48 67 47
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_0
timestamp 1763476864
transform -1 0 1476 0 1 3151
box -96 -124 67 124
use M1_POLY2$$45109292_512x8m81  M1_POLY2$$45109292_512x8m81_0
timestamp 1763476864
transform 1 0 2073 0 1 3335
box -289 -48 289 48
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1763476864
transform 1 0 2475 0 1 498
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1763476864
transform 1 0 2961 0 1 469
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_2
timestamp 1763476864
transform 1 0 2348 0 1 1698
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_3
timestamp 1763476864
transform 1 0 2527 0 1 1826
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_4
timestamp 1763476864
transform 1 0 1824 0 1 498
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_5
timestamp 1763476864
transform 1 0 1986 0 1 498
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_6
timestamp 1763476864
transform 1 0 2331 0 1 498
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_7
timestamp 1763476864
transform 1 0 1459 0 1 541
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_8
timestamp 1763476864
transform 1 0 942 0 1 499
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_9
timestamp 1763476864
transform 1 0 1568 0 1 1687
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_10
timestamp 1763476864
transform 1 0 1317 0 1 541
box -36 -36 36 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_0
timestamp 1763476864
transform 1 0 2019 0 1 2635
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_1
timestamp 1763476864
transform 1 0 1671 0 1 1866
box -62 -36 62 36
use M1_PSUB$$44997676_512x8m81  M1_PSUB$$44997676_512x8m81_0
timestamp 1763476864
transform 1 0 3357 0 -1 1460
box -165 -114 166 114
use M1_PSUB$$44997676_512x8m81  M1_PSUB$$44997676_512x8m81_1
timestamp 1763476864
transform 1 0 -106 0 -1 1460
box -165 -114 166 114
use M1_PSUB_285_512x8m81  M1_PSUB_285_512x8m81_0
timestamp 1763476864
transform 1 0 3413 0 -1 745
box -118 -58 111 57
use M1_PSUB_285_512x8m81  M1_PSUB_285_512x8m81_1
timestamp 1763476864
transform 1 0 -171 0 -1 745
box -118 -58 111 57
use M2_M1$$43374636_512x8m81  M2_M1$$43374636_512x8m81_0
timestamp 1763476864
transform 1 0 170 0 1 1003
box -119 -123 119 123
use M2_M1$$45002796_512x8m81  M2_M1$$45002796_512x8m81_0
timestamp 1763476864
transform 1 0 2144 0 1 926
box -783 -46 783 46
use M2_M1$$45003820_512x8m81  M2_M1$$45003820_512x8m81_0
timestamp 1763476864
transform 1 0 3320 0 1 1079
box -119 -198 119 198
use M2_M1c$$203396140_512x8m81  M2_M1c$$203396140_512x8m81_0
timestamp 1763476864
transform 1 0 697 0 1 2781
box -108 -46 108 46
use M3_M2$$45005868_512x8m81  M3_M2$$45005868_512x8m81_0
timestamp 1763476864
transform 1 0 2144 0 1 926
box -783 -46 783 46
use M3_M2$$45006892_512x8m81  M3_M2$$45006892_512x8m81_0
timestamp 1763476864
transform 1 0 3320 0 1 1079
box -119 -198 119 198
use M3_M2$$45008940_512x8m81  M3_M2$$45008940_512x8m81_0
timestamp 1763476864
transform 1 0 170 0 1 1003
box -119 -123 119 123
use nmos_1p2$$45100076_512x8m81  nmos_1p2$$45100076_512x8m81_0
timestamp 1763476864
transform -1 0 2814 0 -1 1610
box -130 -44 263 287
use nmos_1p2$$45101100_512x8m81  nmos_1p2$$45101100_512x8m81_0
timestamp 1763476864
transform 1 0 241 0 1 598
box -214 -44 660 150
use nmos_1p2$$45102124_512x8m81  nmos_1p2$$45102124_512x8m81_0
timestamp 1763476864
transform -1 0 1106 0 -1 1610
box -270 -44 928 255
use nmos_1p2$$45103148_512x8m81  nmos_1p2$$45103148_512x8m81_0
timestamp 1763476864
transform -1 0 2233 0 -1 1610
box -242 -44 792 310
use nmos_5p04310591302012_512x8m81  nmos_5p04310591302012_512x8m81_0
timestamp 1763476864
transform -1 0 3188 0 1 3504
box -171 -44 541 255
use nmos_5p04310591302023_512x8m81  nmos_5p04310591302023_512x8m81_0
timestamp 1763476864
transform 1 0 2185 0 1 618
box -124 -44 285 100
use nmos_5p04310591302023_512x8m81  nmos_5p04310591302023_512x8m81_1
timestamp 1763476864
transform 1 0 1181 0 1 618
box -124 -44 285 100
use nmos_5p04310591302023_512x8m81  nmos_5p04310591302023_512x8m81_2
timestamp 1763476864
transform 1 0 1688 0 1 618
box -124 -44 285 100
use nmos_5p04310591302028_512x8m81  nmos_5p04310591302028_512x8m81_0
timestamp 1763476864
transform 1 0 849 0 1 3504
box -184 -44 692 255
use nmos_5p04310591302028_512x8m81  nmos_5p04310591302028_512x8m81_1
timestamp 1763476864
transform 1 0 1838 0 1 3504
box -184 -44 692 255
use nmos_5p04310591302032_512x8m81  nmos_5p04310591302032_512x8m81_0
timestamp 1763476864
transform -1 0 304 0 1 3656
box -116 -44 277 150
use nmos_5p04310591302033_512x8m81  nmos_5p04310591302033_512x8m81_0
timestamp 1763476864
transform 1 0 2653 0 1 618
box -92 -44 148 100
use nmos_5p04310591302034_512x8m81  nmos_5p04310591302034_512x8m81_0
timestamp 1763476864
transform 1 0 2985 0 1 572
box -88 -44 144 178
use pmos_1p2$$45095980_512x8m81  pmos_1p2$$45095980_512x8m81_0
timestamp 1763476864
transform -1 0 3017 0 1 2863
box -440 -86 1408 339
use pmos_1p2$$46281772_512x8m81  pmos_1p2$$46281772_512x8m81_0
timestamp 1763476864
transform -1 0 2943 0 -1 2555
box -244 -86 481 509
use pmos_1p2$$46281772_512x8m81  pmos_1p2$$46281772_512x8m81_1
timestamp 1763476864
transform -1 0 2317 0 -1 2555
box -244 -86 481 509
use pmos_1p2$$46282796_512x8m81  pmos_1p2$$46282796_512x8m81_0
timestamp 1763476864
transform 1 0 256 0 1 82
box -300 -86 746 297
use pmos_1p2$$46283820_512x8m81  pmos_1p2$$46283820_512x8m81_0
timestamp 1763476864
transform -1 0 1323 0 -1 2540
box -440 -86 1408 467
use pmos_1p2$$46284844_512x8m81  pmos_1p2$$46284844_512x8m81_0
timestamp 1763476864
transform 1 0 3027 0 1 137
box -216 -86 348 245
use pmos_1p2$$46285868_512x8m81  pmos_1p2$$46285868_512x8m81_0
timestamp 1763476864
transform 1 0 1248 0 1 2938
box -188 -86 216 297
use pmos_1p2$$46286892_512x8m81  pmos_1p2$$46286892_512x8m81_0
timestamp 1763476864
transform 1 0 823 0 1 2938
box -244 -86 481 297
use pmos_1p2$$46287916_512x8m81  pmos_1p2$$46287916_512x8m81_0
timestamp 1763476864
transform -1 0 290 0 1 2932
box -216 -86 348 404
use pmos_5p04310591302027_512x8m81  pmos_5p04310591302027_512x8m81_0
timestamp 1763476864
transform 1 0 2185 0 1 207
box -202 -86 362 198
use pmos_5p04310591302027_512x8m81  pmos_5p04310591302027_512x8m81_1
timestamp 1763476864
transform 1 0 1181 0 1 207
box -202 -86 362 198
use pmos_5p04310591302027_512x8m81  pmos_5p04310591302027_512x8m81_2
timestamp 1763476864
transform 1 0 1688 0 1 207
box -202 -86 362 198
use pmos_5p04310591302038_512x8m81  pmos_5p04310591302038_512x8m81_0
timestamp 1763476864
transform 1 0 2653 0 1 233
box -174 -86 230 198
use po_m1_512x8m81  po_m1_512x8m81_0
timestamp 1763476864
transform 1 0 1920 0 1 1008
box -21 0 113 95
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_0
timestamp 1763476864
transform 1 0 2232 0 1 88
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_1
timestamp 1763476864
transform 1 0 1726 0 1 88
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_2
timestamp 1763476864
transform -1 0 2465 0 -1 1575
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_3
timestamp 1763476864
transform 1 0 3436 0 1 581
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_4
timestamp 1763476864
transform 1 0 3436 0 1 1353
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_5
timestamp 1763476864
transform 1 0 3220 0 1 88
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_6
timestamp 1763476864
transform 1 0 2903 0 1 88
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_7
timestamp 1763476864
transform 1 0 2759 0 1 88
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_8
timestamp 1763476864
transform -1 0 2933 0 -1 1575
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_9
timestamp 1763476864
transform -1 0 2620 0 -1 1575
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_10
timestamp 1763476864
transform -1 0 1521 0 -1 1575
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_11
timestamp 1763476864
transform 1 0 50 0 1 135
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_12
timestamp 1763476864
transform -1 0 -184 0 -1 388
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_13
timestamp 1763476864
transform -1 0 1054 0 -1 1575
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_14
timestamp 1763476864
transform 1 0 -249 0 1 581
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_15
timestamp 1763476864
transform 1 0 -249 0 1 1353
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_16
timestamp 1763476864
transform 1 0 1218 0 1 88
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_17
timestamp 1763476864
transform 1 0 677 0 1 133
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_18
timestamp 1763476864
transform 1 0 364 0 1 134
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_19
timestamp 1763476864
transform 1 0 -249 0 1 2174
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_20
timestamp 1763476864
transform -1 0 79 0 -1 3871
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_21
timestamp 1763476864
transform -1 0 84 0 -1 3086
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_22
timestamp 1763476864
transform -1 0 745 0 -1 3811
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_23
timestamp 1763476864
transform -1 0 1052 0 -1 3811
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_24
timestamp 1763476864
transform -1 0 1379 0 -1 3811
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_25
timestamp 1763476864
transform -1 0 420 0 -1 3871
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_26
timestamp 1763476864
transform -1 0 408 0 -1 3086
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_27
timestamp 1763476864
transform -1 0 746 0 -1 3116
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_28
timestamp 1763476864
transform -1 0 1054 0 -1 3086
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_29
timestamp 1763476864
transform -1 0 83 0 -1 2545
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_30
timestamp 1763476864
transform -1 0 1054 0 -1 2545
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_31
timestamp 1763476864
transform -1 0 -184 0 -1 3885
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_32
timestamp 1763476864
transform -1 0 1359 0 -1 3086
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_33
timestamp 1763476864
transform 1 0 -249 0 1 2578
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_34
timestamp 1763476864
transform 1 0 3436 0 1 2174
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_35
timestamp 1763476864
transform 1 0 3436 0 1 2501
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_36
timestamp 1763476864
transform -1 0 2619 0 -1 2502
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_37
timestamp 1763476864
transform -1 0 2934 0 -1 2502
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_38
timestamp 1763476864
transform -1 0 2308 0 -1 2502
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_39
timestamp 1763476864
transform -1 0 2007 0 -1 2502
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_40
timestamp 1763476864
transform -1 0 1789 0 -1 3103
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_41
timestamp 1763476864
transform -1 0 2095 0 -1 3103
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_42
timestamp 1763476864
transform -1 0 2404 0 -1 3103
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_43
timestamp 1763476864
transform -1 0 2722 0 -1 3103
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_44
timestamp 1763476864
transform -1 0 3034 0 -1 3103
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_45
timestamp 1763476864
transform -1 0 3348 0 -1 3103
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_46
timestamp 1763476864
transform -1 0 2720 0 -1 3811
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_47
timestamp 1763476864
transform -1 0 3033 0 -1 3811
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_48
timestamp 1763476864
transform -1 0 3349 0 -1 3811
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_49
timestamp 1763476864
transform -1 0 3092 0 -1 2074
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_50
timestamp 1763476864
transform -1 0 2777 0 -1 2074
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_51
timestamp 1763476864
transform -1 0 1672 0 -1 2515
box -9 0 73 215
use via1_R90_512x8m81  via1_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 1695 1 0 1852
box 0 0 65 89
use via1_x2_512x8m81  via1_x2_512x8m81_0
timestamp 1763476864
transform 1 0 1736 0 1 590
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_1
timestamp 1763476864
transform 1 0 2242 0 1 590
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_2
timestamp 1763476864
transform 1 0 2750 0 1 590
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_3
timestamp 1763476864
transform 1 0 2907 0 1 590
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_4
timestamp 1763476864
transform 1 0 3063 0 1 542
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_5
timestamp 1763476864
transform 1 0 1052 0 1 355
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_6
timestamp 1763476864
transform 1 0 1274 0 1 590
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_7
timestamp 1763476864
transform 1 0 50 0 1 590
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_8
timestamp 1763476864
transform 1 0 344 0 1 590
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_9
timestamp 1763476864
transform 1 0 674 0 1 590
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_10
timestamp 1763476864
transform -1 0 1501 0 -1 3231
box -8 0 72 222
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 3128 1 0 1058
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_1
timestamp 1763476864
transform 0 -1 3000 1 0 434
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_2
timestamp 1763476864
transform 0 -1 817 1 0 1058
box -8 0 72 215
use via1_x2_R270_512x8m81  via1_x2_R270_512x8m81_0
timestamp 1763476864
transform 0 1 2158 -1 0 1734
box -8 0 75 215
use via1_x2_R270_512x8m81  via1_x2_R270_512x8m81_1
timestamp 1763476864
transform 0 1 994 -1 0 807
box -8 0 75 215
use via1_x2_R270_512x8m81  via1_x2_R270_512x8m81_2
timestamp 1763476864
transform 0 1 1944 -1 0 2676
box -8 0 75 215
use via1_x2_R270_512x8m81  via1_x2_R270_512x8m81_3
timestamp 1763476864
transform 0 1 1526 -1 0 1731
box -8 0 75 215
use via1_x2_R270_512x8m81  via1_x2_R270_512x8m81_4
timestamp 1763476864
transform 0 1 1592 -1 0 3383
box -8 0 75 215
use via2_x2_512x8m81  via2_x2_512x8m81_0
timestamp 1763476864
transform 1 0 2242 0 1 582
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_1
timestamp 1763476864
transform 1 0 1736 0 1 582
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_2
timestamp 1763476864
transform 1 0 2750 0 1 582
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_3
timestamp 1763476864
transform 1 0 2907 0 1 582
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_4
timestamp 1763476864
transform 1 0 674 0 1 582
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_5
timestamp 1763476864
transform 1 0 344 0 1 582
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_6
timestamp 1763476864
transform 1 0 50 0 1 582
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_7
timestamp 1763476864
transform 1 0 1274 0 1 582
box -9 0 74 222
use via2_x2_R90_512x8m81  via2_x2_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 1747 1 0 1860
box -9 0 73 215
<< labels >>
rlabel metal3 s 1678 2661 1678 2661 4 vdd
port 1 nsew
rlabel metal3 s 1514 3810 1514 3810 4 vss
port 2 nsew
rlabel metal3 s 1601 742 1601 742 4 vss
port 2 nsew
rlabel metal3 s 173 1005 173 1005 4 men
port 3 nsew
rlabel metal3 s 1601 1505 1601 1505 4 vss
port 2 nsew
rlabel metal3 s 1042 265 1042 265 4 vdd
port 1 nsew
rlabel metal1 s 1019 1808 1019 1808 4 pcb
port 4 nsew
rlabel metal1 s 2846 3895 2846 3895 4 se
port 5 nsew
<< properties >>
string path 20.320 27.120 20.320 27.785 22.565 27.785 22.565 26.905 
<< end >>
