magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< nsubdiff >>
rect -53 80 53 113
rect -53 -80 -23 80
rect 23 -80 53 80
rect -53 -112 53 -80
<< nsubdiffcont >>
rect -23 -80 23 80
<< metal1 >>
rect -40 80 40 99
rect -40 -80 -23 80
rect 23 -80 40 80
rect -40 -99 40 -80
<< end >>
