magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< nwell >>
rect -202 -86 362 1264
<< pmos >>
rect -28 0 28 1178
rect 132 0 188 1178
<< pdiff >>
rect -116 1165 -28 1178
rect -116 14 -103 1165
rect -57 14 -28 1165
rect -116 0 -28 14
rect 28 1165 132 1178
rect 28 14 57 1165
rect 103 14 132 1165
rect 28 0 132 14
rect 188 1165 276 1178
rect 188 14 217 1165
rect 263 14 276 1165
rect 188 0 276 14
<< pdiffc >>
rect -103 14 -57 1165
rect 57 14 103 1165
rect 217 14 263 1165
<< polysilicon >>
rect -28 1178 28 1222
rect 132 1178 188 1222
rect -28 -44 28 0
rect 132 -44 188 0
<< metal1 >>
rect -103 1165 -57 1178
rect -103 0 -57 14
rect 57 1165 103 1178
rect 57 0 103 14
rect 217 1165 263 1178
rect 217 0 263 14
<< labels >>
flabel pdiffc 80 589 80 589 0 FreeSans 186 0 0 0 D
flabel pdiffc -68 589 -68 589 0 FreeSans 186 0 0 0 S
flabel pdiffc 228 589 228 589 0 FreeSans 186 0 0 0 S
<< end >>
