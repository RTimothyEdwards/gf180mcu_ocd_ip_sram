magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -119 324 119 351
rect -119 -124 -93 324
rect 93 -124 119 324
rect -119 -151 119 -124
<< via2 >>
rect -93 -124 93 324
<< metal3 >>
rect -119 324 119 351
rect -119 -124 -93 324
rect 93 -124 119 324
rect -119 -151 119 -124
<< end >>
