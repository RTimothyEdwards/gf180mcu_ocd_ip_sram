magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< psubdiff >>
rect -91 23 91 56
rect -91 -23 -23 23
rect 23 -23 91 23
rect -91 -56 91 -23
<< psubdiffcont >>
rect -23 -23 23 23
<< metal1 >>
rect -40 23 40 42
rect -40 -23 -23 23
rect 23 -23 40 23
rect -40 -42 40 -23
<< end >>
