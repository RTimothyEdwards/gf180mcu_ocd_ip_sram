magic
tech gf180mcuD
magscale 1 10
timestamp 1765921700
<< error_s >>
rect 1572 13654 1611 13655
rect 1645 13654 1684 13655
rect 1770 13654 1809 13655
rect 1843 13654 1882 13655
rect 1968 13654 2007 13655
rect 2041 13654 2080 13655
rect 2852 13654 2891 13655
rect 2925 13654 2964 13655
rect 3050 13654 3089 13655
rect 3123 13654 3162 13655
rect 3248 13654 3287 13655
rect 3321 13654 3360 13655
rect 6737 13654 6776 13655
rect 6810 13654 6849 13655
rect 6935 13654 6974 13655
rect 7008 13654 7047 13655
rect 7133 13654 7172 13655
rect 7206 13654 7245 13655
rect 8017 13654 8056 13655
rect 8090 13654 8129 13655
rect 8215 13654 8254 13655
rect 8288 13654 8327 13655
rect 8413 13654 8452 13655
rect 8486 13654 8525 13655
<< nwell >>
rect 17442 18870 18301 19318
rect 17262 8699 17293 8720
rect 18106 8699 18193 8720
rect 18983 8699 19055 8720
rect 14494 7349 15036 7710
rect 16382 7653 19055 8699
rect 14517 6396 14632 6429
rect 17262 5806 17293 7653
rect 18106 5377 18193 7653
rect 18983 5471 19055 7653
rect 5846 2204 6015 2612
<< metal1 >>
rect 282 19904 375 19938
rect 282 19700 303 19904
rect 355 19700 375 19904
rect 1143 19797 1270 19844
rect 282 2508 375 19700
rect 4808 13607 4899 13808
rect 535 13513 4899 13607
rect 535 9206 625 13513
rect 6001 13448 6092 13799
rect 704 13354 6092 13448
rect 704 9470 795 13354
rect 9952 13289 10042 13787
rect 873 13196 10042 13289
rect 11136 13333 11226 13841
rect 17292 13492 17383 13878
rect 18476 13651 18566 13878
rect 19660 13809 19753 13878
rect 19660 13716 20202 13809
rect 19660 13715 19753 13716
rect 18476 13557 20033 13651
rect 17292 13399 19864 13492
rect 11136 13240 19695 13333
rect 873 9675 963 13196
rect 873 9586 1290 9675
rect 704 9361 1121 9470
rect 535 9099 952 9206
rect 861 2264 952 9099
rect 1031 2264 1121 9361
rect 1199 2264 1290 9586
rect 14693 8441 14743 8570
rect 15017 8441 15068 8575
rect 15336 8441 15386 8561
rect 14693 8391 15386 8441
rect 14710 8390 15369 8391
rect 15701 2862 15748 2864
rect 14532 2813 15748 2862
rect 9200 1985 10308 2033
rect 15701 2007 15748 2813
rect 19604 2121 19695 13240
rect 19773 2121 19864 13399
rect 19943 2121 20033 13557
rect 20111 2121 20202 13716
rect 20664 2508 20757 19906
rect 282 1612 6454 1931
rect 9200 648 9248 1985
rect 19488 1612 20590 1931
<< metal2 >>
rect 451 2667 1043 20627
rect 12009 19735 12100 19828
rect 12255 19735 12345 19828
rect 13153 19735 13244 19828
rect 13402 19735 13492 19828
rect 14298 19735 14389 19828
rect 14538 19735 14628 19828
rect 15439 19735 15529 19828
rect 15691 19735 15781 19828
rect 1635 19576 1725 19670
rect 1883 19576 1974 19670
rect 2887 19576 2978 19670
rect 3141 19576 3231 19670
rect 6799 19576 6890 19670
rect 7049 19576 7139 19670
rect 8052 19576 8143 19670
rect 8306 19576 8397 19670
rect 282 702 375 2509
rect 451 1612 760 2667
rect 861 702 952 2509
rect 1031 702 1121 2509
rect 1199 702 1290 2509
rect 2359 702 2452 3052
rect 3542 702 3636 3068
rect 4727 702 4821 3059
rect 6274 2924 6364 3076
rect 5693 2830 6364 2924
rect 11423 2855 11480 2857
rect 5693 1008 5783 2830
rect 11353 2816 11480 2855
rect 6216 1816 6454 2724
rect 11423 744 11480 2816
rect 15128 1600 15375 4119
rect 19972 2667 20588 20627
rect 15998 702 16092 2132
rect 19604 702 19695 2519
rect 19773 702 19864 2519
rect 19943 702 20033 2519
rect 20111 702 20202 2519
rect 20279 1612 20588 2667
rect 20664 820 20757 2509
<< metal3 >>
rect 451 19991 20588 20627
rect 282 19864 20757 19906
rect 282 19690 20667 19864
rect 20753 19690 20757 19864
rect 11520 14633 11610 15111
rect 16190 14633 16350 15110
rect 16290 14186 16360 14552
rect 19677 12097 19767 12190
rect 19677 11859 19767 11952
rect 19677 11621 19767 11714
rect 19677 11383 19767 11476
rect 19677 11145 19767 11238
rect 19677 10907 19767 11000
rect 19677 10668 19767 10762
rect 19677 10430 19767 10524
use gen_3v1024x8_3v1024x8m81  gen_3v1024x8_3v1024x8m81_0
timestamp 1765921700
transform 1 0 9916 0 1 2199
box -12453 -1374 12336 10979
use M1_NACTIVE4310591302047_3v1024x8m81  M1_NACTIVE4310591302047_3v1024x8m81_0
timestamp 1764525316
transform 0 -1 18221 1 0 19090
box -96 -86 96 86
use M1_NACTIVE4310591302047_3v1024x8m81  M1_NACTIVE4310591302047_3v1024x8m81_1
timestamp 1764525316
transform 0 -1 17500 1 0 19099
box -96 -86 96 86
use M1_PACTIVE4310591302048_3v1024x8m81  M1_PACTIVE4310591302048_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2440 0 1 19821
box -1152 -36 1153 36
use M1_PACTIVE4310591302048_3v1024x8m81  M1_PACTIVE4310591302048_3v1024x8m81_1
timestamp 1764525316
transform 1 0 7592 0 1 19821
box -1152 -36 1153 36
use M1_PACTIVE4310591302049_3v1024x8m81  M1_PACTIVE4310591302049_3v1024x8m81_0
timestamp 1764525316
transform 1 0 16713 0 1 19808
box -457 -36 457 36
use M2_M1$$43375660_3v1024x8m81  M2_M1$$43375660_3v1024x8m81_0
timestamp 1764525316
transform -1 0 20710 0 1 19812
box -43 -122 43 122
use M2_M1$$43375660_3v1024x8m81  M2_M1$$43375660_3v1024x8m81_1
timestamp 1764525316
transform -1 0 20710 0 1 2387
box -43 -122 43 122
use M2_M1$$43375660_3v1024x8m81  M2_M1$$43375660_3v1024x8m81_2
timestamp 1764525316
transform 1 0 329 0 1 19802
box -43 -122 43 122
use M2_M1$$43375660_3v1024x8m81  M2_M1$$43375660_3v1024x8m81_3
timestamp 1764525316
transform 1 0 329 0 1 2387
box -43 -122 43 122
use M2_M1$$199746604_3v1024x8m81  M2_M1$$199746604_3v1024x8m81_0
timestamp 1764525316
transform 1 0 605 0 1 1771
box -119 -123 119 123
use M2_M1$$199746604_3v1024x8m81  M2_M1$$199746604_3v1024x8m81_1
timestamp 1764525316
transform 1 0 20433 0 1 1771
box -119 -123 119 123
use M2_M1$$199746604_3v1024x8m81  M2_M1$$199746604_3v1024x8m81_2
timestamp 1764525316
transform 1 0 6335 0 1 1697
box -119 -123 119 123
use M2_M1$$201262124_3v1024x8m81  M2_M1$$201262124_3v1024x8m81_0
timestamp 1764525316
transform 1 0 6335 0 1 1884
box -119 -46 119 46
use M2_M1$$202405932_3v1024x8m81  M2_M1$$202405932_3v1024x8m81_0
timestamp 1764525316
transform 1 0 20157 0 1 2320
box -44 -198 44 198
use M2_M1$$202405932_3v1024x8m81  M2_M1$$202405932_3v1024x8m81_1
timestamp 1764525316
transform 1 0 19988 0 1 2320
box -44 -198 44 198
use M2_M1$$202405932_3v1024x8m81  M2_M1$$202405932_3v1024x8m81_2
timestamp 1764525316
transform 1 0 19819 0 1 2320
box -44 -198 44 198
use M2_M1$$202405932_3v1024x8m81  M2_M1$$202405932_3v1024x8m81_3
timestamp 1764525316
transform 1 0 19649 0 1 2320
box -44 -198 44 198
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1245 0 1 2387
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_1
timestamp 1764525316
transform 1 0 1075 0 1 2387
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_2
timestamp 1764525316
transform 1 0 907 0 1 2387
box -45 -122 45 123
use M3_M2$$43368492_3v1024x8m81  M3_M2$$43368492_3v1024x8m81_0
timestamp 1764525316
transform -1 0 20710 0 1 19812
box -44 -123 44 123
use M3_M2$$43368492_3v1024x8m81  M3_M2$$43368492_3v1024x8m81_1
timestamp 1764525316
transform 1 0 329 0 1 19812
box -44 -123 44 123
use M3_M2$$201255980_3v1024x8m81  M3_M2$$201255980_3v1024x8m81_0
timestamp 1764525316
transform -1 0 20640 0 1 1028
box -119 -46 119 46
use M3_M2$$201255980_3v1024x8m81  M3_M2$$201255980_3v1024x8m81_1
timestamp 1764525316
transform 1 0 399 0 1 1028
box -119 -46 119 46
use M3_M2$$201255980_3v1024x8m81  M3_M2$$201255980_3v1024x8m81_2
timestamp 1764525316
transform 1 0 5738 0 1 1028
box -119 -46 119 46
use M3_M2$$201401388_3v1024x8m81  M3_M2$$201401388_3v1024x8m81_0
timestamp 1764525316
transform 1 0 20280 0 1 20309
box -266 -275 266 275
use M3_M2$$201401388_3v1024x8m81  M3_M2$$201401388_3v1024x8m81_1
timestamp 1764525316
transform 1 0 759 0 1 20309
box -266 -275 266 275
use M3_M2$$201401388_3v1024x8m81  M3_M2$$201401388_3v1024x8m81_2
timestamp 1764525316
transform 1 0 20280 0 1 8482
box -266 -275 266 275
use M3_M24310591302050_3v1024x8m81  M3_M24310591302050_3v1024x8m81_0
timestamp 1764525316
transform 1 0 15254 0 1 1756
box -99 -99 99 99
use M3_M24310591302050_3v1024x8m81  M3_M24310591302050_3v1024x8m81_1
timestamp 1764525316
transform 1 0 15254 0 1 2372
box -99 -99 99 99
use prexdec_top_3v1024x8m81  prexdec_top_3v1024x8m81_0
timestamp 1765921700
transform 1 0 949 0 1 11846
box 21 1806 19120 8780
use ypredec1_3v1024x8m81  ypredec1_3v1024x8m81_0
timestamp 1765921204
transform 1 0 1092 0 1 2092
box 125 53 18674 11111
<< labels >>
flabel metal1 s 9219 762 9219 762 0 FreeSans 700 0 0 0 GWEN
port 51 nsew
flabel metal1 s 15717 2437 15717 2437 0 FreeSans 700 0 0 0 GWE
port 50 nsew
rlabel metal2 s 1075 748 1075 748 4 A[8]
port 49 nsew
rlabel metal2 s 19819 748 19819 748 4 A[5]
port 48 nsew
rlabel metal2 s 19988 748 19988 748 4 A[4]
port 47 nsew
rlabel metal2 s 20157 748 20157 748 4 A[3]
port 46 nsew
rlabel metal2 s 19649 748 19649 748 4 A[6]
port 45 nsew
rlabel metal2 s 3589 748 3589 748 4 A[1]
port 44 nsew
rlabel metal2 s 2405 748 2405 748 4 A[2]
port 43 nsew
rlabel metal2 s 329 748 329 748 4 CLK
port 42 nsew
rlabel metal2 s 1245 748 1245 748 4 A[7]
port 41 nsew
rlabel metal2 s 907 748 907 748 4 A[9]
port 40 nsew
rlabel metal2 s 16046 748 16046 748 4 CEN
port 32 nsew
rlabel metal2 s 4774 748 4774 748 4 A[0]
port 31 nsew
flabel metal2 s 11449 762 11449 762 0 FreeSans 700 0 0 0 IGWEN
port 21 nsew
flabel metal3 s 4365 6277 4365 6277 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 4365 3413 4365 3413 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 5796 2441 5796 2441 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 4365 4149 4365 4149 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 4365 8014 4365 8014 0 FreeSans 313 0 0 0 VSS
port 1 nsew
rlabel metal3 s 19569 5213 19569 5213 4 tblhl
port 20 nsew
rlabel metal3 s 19722 12144 19722 12144 4 RYS[7]
port 3 nsew
rlabel metal3 s 19722 11905 19722 11905 4 RYS[6]
port 4 nsew
rlabel metal3 s 19722 11667 19722 11667 4 RYS[5]
port 5 nsew
rlabel metal3 s 19722 11429 19722 11429 4 RYS[4]
port 6 nsew
rlabel metal3 s 19722 11191 19722 11191 4 RYS[3]
port 7 nsew
rlabel metal3 s 19722 10953 19722 10953 4 RYS[2]
port 8 nsew
rlabel metal3 s 19722 10715 19722 10715 4 RYS[1]
port 9 nsew
rlabel metal3 s 19722 10477 19722 10477 4 RYS[0]
port 10 nsew
flabel metal3 s 5488 1266 5488 1266 0 FreeSans 313 0 0 0 VSS
port 1 nsew
rlabel metal3 s 18802 20309 18802 20309 4 men
port 18 nsew
flabel metal3 s 5295 2946 5295 2946 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 6656 1754 6656 1754 0 FreeSans 313 0 0 0 VDD
port 2 nsew
rlabel metal2 s 15484 19781 15484 19781 4 xa[1]
port 39 nsew
rlabel metal2 s 15736 19781 15736 19781 4 xa[0]
port 38 nsew
rlabel metal2 s 14583 19781 14583 19781 4 xa[2]
port 30 nsew
rlabel metal2 s 14343 19781 14343 19781 4 xa[3]
port 29 nsew
rlabel metal2 s 13447 19781 13447 19781 4 xa[4]
port 28 nsew
rlabel metal2 s 13198 19781 13198 19781 4 xa[5]
port 27 nsew
rlabel metal2 s 12300 19781 12300 19781 4 xa[6]
port 26 nsew
rlabel metal2 s 12054 19781 12054 19781 4 xa[7]
port 25 nsew
rlabel metal2 s 6845 19623 6845 19623 4 xb[3]
port 22 nsew
rlabel metal2 s 8098 19620 8098 19620 4 xb[1]
port 33 nsew
rlabel metal2 s 8351 19620 8351 19620 4 xb[0]
port 24 nsew
rlabel metal2 s 7094 19623 7094 19623 4 xb[2]
port 23 nsew
rlabel metal2 s 8068 19628 8068 19628 4 xb[1]
port 33 nsew
rlabel metal2 s 8376 19641 8376 19641 4 xb[0]
port 24 nsew
rlabel metal2 s 7114 19658 7114 19658 4 xb[2]
port 23 nsew
rlabel metal2 s 6808 19653 6808 19653 4 xb[3]
port 22 nsew
rlabel metal2 s 3186 19620 3186 19620 4 xc[0]
port 37 nsew
rlabel metal2 s 1929 19623 1929 19623 4 xc[2]
port 36 nsew
rlabel metal2 s 2933 19620 2933 19620 4 xc[1]
port 35 nsew
rlabel metal2 s 1680 19623 1680 19623 4 xc[3]
port 34 nsew
rlabel metal3 s 1263 10467 1263 10467 4 LYS[0]
port 11 nsew
rlabel metal3 s 1263 10705 1263 10705 4 LYS[1]
port 12 nsew
rlabel metal3 s 1263 10943 1263 10943 4 LYS[2]
port 13 nsew
rlabel metal3 s 1263 11181 1263 11181 4 LYS[3]
port 14 nsew
rlabel metal3 s 1263 11895 1263 11895 4 LYS[6]
port 15 nsew
rlabel metal3 s 1263 11657 1263 11657 4 LYS[5]
port 16 nsew
rlabel metal3 s 1263 11419 1263 11419 4 LYS[4]
port 17 nsew
rlabel metal3 s 1263 12134 1263 12134 4 LYS[7]
port 19 nsew
flabel metal3 s 4385 12709 4385 12709 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 3755 14336 3755 14336 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 3755 14822 3755 14822 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 3775 13901 3775 13901 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 4355 19382 4355 19382 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 4115 18708 4115 18708 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 4005 18116 4005 18116 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 3945 16834 3945 16834 0 FreeSans 313 0 0 0 VDD
port 2 nsew
<< properties >>
string path 81.095 8.115 81.735 8.115 81.735 -9.165 
<< end >>
