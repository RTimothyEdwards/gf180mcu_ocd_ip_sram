magic
tech gf180mcuD
magscale 1 10
timestamp 1765833244
<< psubdiff >>
rect -522 23 522 36
rect -522 -23 -509 23
rect 509 -23 522 23
rect -522 -36 522 -23
<< psubdiffcont >>
rect -509 -23 509 23
<< metal1 >>
rect -517 23 517 30
rect -517 -23 -509 23
rect 509 -23 517 23
rect -517 -30 517 -23
<< end >>
