magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nwell >>
rect -174 -86 230 701
<< pmos >>
rect 0 0 56 615
<< pdiff >>
rect -88 602 0 615
rect -88 13 -75 602
rect -29 13 0 602
rect -88 0 0 13
rect 56 602 144 615
rect 56 13 85 602
rect 131 13 144 602
rect 56 0 144 13
<< pdiffc >>
rect -75 13 -29 602
rect 85 13 131 602
<< polysilicon >>
rect 0 615 56 659
rect 0 -44 56 0
<< metal1 >>
rect -75 602 -29 615
rect -75 0 -29 13
rect 85 602 131 615
rect 85 0 131 13
<< labels >>
flabel pdiffc -40 307 -40 307 0 FreeSans 186 0 0 0 S
flabel pdiffc 96 307 96 307 0 FreeSans 186 0 0 0 D
<< end >>
