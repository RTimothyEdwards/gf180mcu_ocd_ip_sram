magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< nwell >>
rect -202 -86 362 1079
<< pmos >>
rect -28 0 28 993
rect 132 0 188 993
<< pdiff >>
rect -116 980 -28 993
rect -116 13 -103 980
rect -57 13 -28 980
rect -116 0 -28 13
rect 28 980 132 993
rect 28 13 57 980
rect 103 13 132 980
rect 28 0 132 13
rect 188 980 276 993
rect 188 13 217 980
rect 263 13 276 980
rect 188 0 276 13
<< pdiffc >>
rect -103 13 -57 980
rect 57 13 103 980
rect 217 13 263 980
<< polysilicon >>
rect -28 993 28 1037
rect 132 993 188 1037
rect -28 -44 28 0
rect 132 -44 188 0
<< metal1 >>
rect -103 980 -57 993
rect -103 0 -57 13
rect 57 980 103 993
rect 57 0 103 13
rect 217 980 263 993
rect 217 0 263 13
<< labels >>
flabel pdiffc 80 496 80 496 0 FreeSans 186 0 0 0 D
flabel pdiffc -68 496 -68 496 0 FreeSans 186 0 0 0 S
flabel pdiffc 228 496 228 496 0 FreeSans 186 0 0 0 S
<< end >>
