magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal2 >>
rect -45 28 635 46
rect -45 -28 -28 28
rect 619 -28 635 28
rect -45 -46 635 -28
<< via2 >>
rect -28 -28 619 28
<< metal3 >>
rect -45 28 635 46
rect -45 -28 -28 28
rect 619 -28 635 28
rect -45 -46 635 -28
<< end >>
