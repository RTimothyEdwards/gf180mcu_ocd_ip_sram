magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -35 527 35 534
rect -35 -527 -28 527
rect 28 -527 35 527
rect -35 -534 35 -527
<< via2 >>
rect -28 -527 28 527
<< metal3 >>
rect -35 527 35 534
rect -35 -527 -28 527
rect 28 -527 35 527
rect -35 -534 35 -527
<< end >>
