magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< nwell >>
rect -202 -86 362 509
<< pmos >>
rect -28 0 28 423
rect 132 0 188 423
<< pdiff >>
rect -116 410 -28 423
rect -116 13 -103 410
rect -57 13 -28 410
rect -116 0 -28 13
rect 28 410 132 423
rect 28 13 57 410
rect 103 13 132 410
rect 28 0 132 13
rect 188 410 276 423
rect 188 13 217 410
rect 263 13 276 410
rect 188 0 276 13
<< pdiffc >>
rect -103 13 -57 410
rect 57 13 103 410
rect 217 13 263 410
<< polysilicon >>
rect -28 423 28 468
rect 132 423 188 468
rect -28 -44 28 0
rect 132 -44 188 0
<< metal1 >>
rect -103 410 -57 423
rect -103 0 -57 13
rect 57 410 103 423
rect 57 0 103 13
rect 217 410 263 423
rect 217 0 263 13
<< labels >>
flabel pdiffc 80 211 80 211 0 FreeSans 186 0 0 0 D
flabel pdiffc -68 211 -68 211 0 FreeSans 186 0 0 0 S
flabel pdiffc 228 211 228 211 0 FreeSans 186 0 0 0 S
<< end >>
