magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< nwell >>
rect 0 4977 984 5167
rect 0 1605 1067 4977
<< polysilicon >>
rect 184 1923 240 2067
rect 488 2004 544 2035
rect 648 2004 704 2035
rect 808 2004 864 2035
rect 488 1945 889 2004
rect 187 1127 243 1617
rect 491 1565 867 1646
rect 491 1127 547 1565
rect 651 1127 707 1565
rect 811 1127 867 1565
<< metal1 >>
rect 109 3936 155 4623
rect 573 3937 619 4624
rect 893 3940 939 4627
rect 183 1616 231 1961
rect 126 1558 231 1616
rect 279 1640 325 2132
rect 573 1827 619 2109
rect 800 1640 846 1966
rect 279 1612 846 1640
rect 279 1593 816 1612
rect 279 1017 325 1593
rect 416 962 464 1435
rect 736 962 784 1435
rect 101 173 182 346
rect 100 0 182 173
rect 571 0 652 346
rect 885 173 966 346
rect 884 0 966 173
<< metal2 >>
rect 428 2248 481 2311
rect 742 2257 795 2319
rect 118 1557 182 1697
rect 428 1425 485 2248
rect 742 1425 800 2257
<< metal3 >>
rect 120 3950 1351 5167
use M1_NWELL4310591302032_256x8m81  M1_NWELL4310591302032_256x8m81_0
timestamp 1763564386
transform 1 0 620 0 1 1838
box -126 -85 127 87
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_0
timestamp 1763564386
transform 1 0 197 0 1 1953
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_1
timestamp 1763564386
transform 1 0 197 0 1 1587
box -36 -36 36 36
use M1_POLY24310591302033_256x8m81  M1_POLY24310591302033_256x8m81_0
timestamp 1763564386
transform 1 0 819 0 1 1974
box -62 -36 62 36
use M1_POLY24310591302033_256x8m81  M1_POLY24310591302033_256x8m81_1
timestamp 1763564386
transform 1 0 789 0 1 1617
box -62 -36 62 36
use M2_M14310591302052_256x8m81  M2_M14310591302052_256x8m81_0
timestamp 1763564386
transform 1 0 611 0 1 4606
box -34 -504 34 504
use M2_M14310591302052_256x8m81  M2_M14310591302052_256x8m81_1
timestamp 1763564386
transform 1 0 925 0 1 4606
box -34 -504 34 504
use M2_M14310591302052_256x8m81  M2_M14310591302052_256x8m81_2
timestamp 1763564386
transform 1 0 141 0 1 4606
box -34 -504 34 504
use M2_M14310591302054_256x8m81  M2_M14310591302054_256x8m81_0
timestamp 1763564386
transform 1 0 768 0 1 1395
box -34 -113 34 113
use M2_M14310591302054_256x8m81  M2_M14310591302054_256x8m81_1
timestamp 1763564386
transform 1 0 455 0 1 1395
box -34 -113 34 113
use M2_M14310591302055_256x8m81  M2_M14310591302055_256x8m81_0
timestamp 1763564386
transform 1 0 152 0 1 1589
box -34 -34 34 34
use M2_M14310591302056_256x8m81  M2_M14310591302056_256x8m81_0
timestamp 1763564386
transform 1 0 768 0 1 3011
box -34 -764 34 764
use M2_M14310591302056_256x8m81  M2_M14310591302056_256x8m81_1
timestamp 1763564386
transform 1 0 455 0 1 3011
box -34 -764 34 764
use M3_M24310591302053_256x8m81  M3_M24310591302053_256x8m81_0
timestamp 1763564386
transform 1 0 141 0 1 4606
box -35 -504 35 504
use M3_M24310591302053_256x8m81  M3_M24310591302053_256x8m81_1
timestamp 1763564386
transform 1 0 925 0 1 4606
box -35 -504 35 504
use M3_M24310591302053_256x8m81  M3_M24310591302053_256x8m81_2
timestamp 1763564386
transform 1 0 611 0 1 4606
box -35 -504 35 504
use nmos_5p04310591302054_256x8m81  nmos_5p04310591302054_256x8m81_0
timestamp 1763564386
transform 1 0 651 0 1 238
box -88 -44 144 891
use nmos_5p04310591302054_256x8m81  nmos_5p04310591302054_256x8m81_1
timestamp 1763564386
transform 1 0 491 0 1 238
box -88 -44 144 891
use nmos_5p04310591302054_256x8m81  nmos_5p04310591302054_256x8m81_2
timestamp 1763564386
transform 1 0 187 0 1 238
box -88 -44 144 891
use nmos_5p04310591302054_256x8m81  nmos_5p04310591302054_256x8m81_3
timestamp 1763564386
transform 1 0 811 0 1 238
box -88 -44 144 891
use pmos_5p04310591302055_256x8m81  pmos_5p04310591302055_256x8m81_0
timestamp 1763564386
transform 1 0 184 0 1 2079
box -174 -86 230 1952
use pmos_5p04310591302055_256x8m81  pmos_5p04310591302055_256x8m81_1
timestamp 1763564386
transform 1 0 488 0 1 2079
box -174 -86 230 1952
use pmos_5p04310591302055_256x8m81  pmos_5p04310591302055_256x8m81_2
timestamp 1763564386
transform 1 0 648 0 1 2079
box -174 -86 230 1952
use pmos_5p04310591302055_256x8m81  pmos_5p04310591302055_256x8m81_3
timestamp 1763564386
transform 1 0 808 0 1 2079
box -174 -86 230 1952
<< properties >>
string path 4.370 15.035 4.370 13.055 
<< end >>
