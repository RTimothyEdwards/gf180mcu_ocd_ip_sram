magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< psubdiff >>
rect -36 114 36 128
rect -36 -114 -23 114
rect 23 -114 36 114
rect -36 -128 36 -114
<< psubdiffcont >>
rect -23 -114 23 114
<< metal1 >>
rect -30 114 30 122
rect -30 -114 -23 114
rect 23 -114 30 114
rect -30 -122 30 -114
<< end >>
