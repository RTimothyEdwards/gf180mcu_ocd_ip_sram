magic
tech gf180mcuD
magscale 1 10
timestamp 1764700137
<< metal1 >>
rect 0 71 67 89
rect 0 18 7 71
rect 59 18 67 71
rect 0 0 67 18
<< via1 >>
rect 7 18 59 71
<< metal2 >>
rect 0 71 67 88
rect 0 18 7 71
rect 59 18 67 71
rect 0 0 67 18
<< end >>
