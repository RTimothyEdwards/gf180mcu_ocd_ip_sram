magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect -174 -86 230 1314
<< pmos >>
rect 0 0 56 1228
<< pdiff >>
rect -88 1215 0 1228
rect -88 13 -75 1215
rect -29 13 0 1215
rect -88 0 0 13
rect 56 1215 144 1228
rect 56 13 85 1215
rect 131 13 144 1215
rect 56 0 144 13
<< pdiffc >>
rect -75 13 -29 1215
rect 85 13 131 1215
<< polysilicon >>
rect 0 1228 56 1272
rect 0 -44 56 0
<< metal1 >>
rect -75 1215 -29 1228
rect -75 0 -29 13
rect 85 1215 131 1228
rect 85 0 131 13
<< labels >>
flabel pdiffc -40 614 -40 614 0 FreeSans 186 0 0 0 S
flabel pdiffc 96 614 96 614 0 FreeSans 186 0 0 0 D
<< end >>
