magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< psubdiff >>
rect -665 23 665 57
rect -665 -23 -632 23
rect 632 -23 665 23
rect -665 -58 665 -23
<< psubdiffcont >>
rect -632 -23 632 23
<< metal1 >>
rect -658 23 658 51
rect -658 -23 -632 23
rect 632 -23 658 23
rect -658 -51 658 -23
<< end >>
