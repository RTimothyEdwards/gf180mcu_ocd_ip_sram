magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< nwell >>
rect -133 -65 160 277
<< polysilicon >>
rect -14 211 41 245
rect -14 -34 41 0
use pmos_5p04310591302014_512x8m81  pmos_5p04310591302014_512x8m81_0
timestamp 1763765945
transform 1 0 -14 0 1 0
box -174 -86 230 297
<< end >>
