* NGSPICE file created from gf180mcu_ocd_ip_sram__sram1024x8m8wm1.ext - technology: gf180mcuD

.subckt pmos_5p0431059130201_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=1.397p pd=7.23u as=1.397p ps=7.23u w=3.175u l=0.28u
.ends

.subckt pmos_1p2$$46889004_3v1024x8m81 pmos_5p0431059130201_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p0431059130201_3v1024x8m81_0/S
Xpmos_5p0431059130201_3v1024x8m81_0 pmos_5p0431059130201_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p0431059130201_3v1024x8m81_0/S pmos_5p0431059130201_3v1024x8m81
.ends

.subckt pmos_5p0431059130206_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.1157p pd=0.965u as=0.1958p ps=1.77u w=0.445u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.1958p pd=1.77u as=0.1157p ps=0.965u w=0.445u l=0.28u
.ends

.subckt pmos_1p2$$46885932_3v1024x8m81 pmos_5p0431059130206_3v1024x8m81_0/D pmos_5p0431059130206_3v1024x8m81_0/S_uq0
+ pmos_5p0431059130206_3v1024x8m81_0/S a_118_89# a_n42_89# w_n133_n65#
Xpmos_5p0431059130206_3v1024x8m81_0 pmos_5p0431059130206_3v1024x8m81_0/D a_n42_89#
+ a_118_89# w_n133_n65# pmos_5p0431059130206_3v1024x8m81_0/S_uq0 pmos_5p0431059130206_3v1024x8m81_0/S
+ pmos_5p0431059130206_3v1024x8m81
.ends

.subckt nmos_5p0431059130207_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=2.794p pd=13.58u as=2.794p ps=13.58u w=6.35u l=0.28u
.ends

.subckt nmos_1p2$$46884908_3v1024x8m81 nmos_5p0431059130207_3v1024x8m81_0/S a_n14_n34#
+ nmos_5p0431059130207_3v1024x8m81_0/D VSUBS
Xnmos_5p0431059130207_3v1024x8m81_0 nmos_5p0431059130207_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p0431059130207_3v1024x8m81_0/S VSUBS nmos_5p0431059130207_3v1024x8m81
.ends

.subckt pmos_5p0431059130209_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.3276p pd=11.46u as=2.3276p ps=11.46u w=5.29u l=0.28u
.ends

.subckt pmos_5p0431059130204_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.794p pd=13.58u as=2.794p ps=13.58u w=6.35u l=0.28u
.ends

.subckt pmos_1p2$$46887980_3v1024x8m81 w_n133_n66# pmos_5p0431059130204_3v1024x8m81_0/S
+ pmos_5p0431059130204_3v1024x8m81_0/D a_n14_n34#
Xpmos_5p0431059130204_3v1024x8m81_0 pmos_5p0431059130204_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p0431059130204_3v1024x8m81_0/S pmos_5p0431059130204_3v1024x8m81
.ends

.subckt pmos_5p0431059130203_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.1378p pd=1.05u as=0.2332p ps=1.94u w=0.53u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.2332p pd=1.94u as=0.1378p ps=1.05u w=0.53u l=0.28u
.ends

.subckt pmos_1p2$$46273580_3v1024x8m81 w_n133_n66# a_n42_n34# pmos_5p0431059130203_3v1024x8m81_0/S
+ a_118_n34# pmos_5p0431059130203_3v1024x8m81_0/D pmos_5p0431059130203_3v1024x8m81_0/S_uq0
Xpmos_5p0431059130203_3v1024x8m81_0 pmos_5p0431059130203_3v1024x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p0431059130203_3v1024x8m81_0/S_uq0 pmos_5p0431059130203_3v1024x8m81_0/S
+ pmos_5p0431059130203_3v1024x8m81
.ends

.subckt nmos_5p04310591302011_3v1024x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.1157p pd=0.965u as=0.1958p ps=1.77u w=0.445u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.1958p pd=1.77u as=0.1157p ps=0.965u w=0.445u l=0.28u
.ends

.subckt nmos_5p0431059130208_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
.ends

.subckt nmos_1p2$$46563372_3v1024x8m81 nmos_5p0431059130208_3v1024x8m81_0/S nmos_5p0431059130208_3v1024x8m81_0/D
+ a_n14_89# VSUBS
Xnmos_5p0431059130208_3v1024x8m81_0 nmos_5p0431059130208_3v1024x8m81_0/D a_n14_89#
+ nmos_5p0431059130208_3v1024x8m81_0/S VSUBS nmos_5p0431059130208_3v1024x8m81
.ends

.subckt nmos_5p04310591302010_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.4642p ps=2.99u w=1.055u l=0.28u
.ends

.subckt nmos_5p0431059130205_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=2.3276p pd=11.46u as=2.3276p ps=11.46u w=5.29u l=0.28u
.ends

.subckt nmos_1p2$$46883884_3v1024x8m81 nmos_5p0431059130205_3v1024x8m81_0/D nmos_5p0431059130205_3v1024x8m81_0/S
+ a_n14_n34# VSUBS
Xnmos_5p0431059130205_3v1024x8m81_0 nmos_5p0431059130205_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p0431059130205_3v1024x8m81_0/S VSUBS nmos_5p0431059130205_3v1024x8m81
.ends

.subckt din_3v1024x8m81 vss datain men db d wep pmos_5p0431059130206_3v1024x8m81_0/D
+ vdd m1_114_5647# VSUBS
Xpmos_1p2$$46889004_3v1024x8m81_0 pmos_1p2$$46889004_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ a_507_5030# vdd d pmos_1p2$$46889004_3v1024x8m81
Xpmos_1p2$$46889004_3v1024x8m81_1 pmos_5p0431059130209_3v1024x8m81_0/S a_507_5030#
+ vdd db pmos_1p2$$46889004_3v1024x8m81
Xpmos_1p2$$46885932_3v1024x8m81_0 nmos_5p04310591302011_3v1024x8m81_1/D nmos_5p04310591302011_3v1024x8m81_1/S_uq0
+ nmos_5p04310591302011_3v1024x8m81_1/S pmos_1p2$$46273580_3v1024x8m81_0/pmos_5p0431059130203_3v1024x8m81_0/D
+ men pmos_5p0431059130206_3v1024x8m81_0/D pmos_1p2$$46885932_3v1024x8m81
Xnmos_1p2$$46884908_3v1024x8m81_0 VSUBS pmos_5p0431059130201_3v1024x8m81_0/S pmos_1p2$$46889004_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ VSUBS nmos_1p2$$46884908_3v1024x8m81
Xpmos_5p0431059130201_3v1024x8m81_0 pmos_5p0431059130206_3v1024x8m81_0/D nmos_5p04310591302011_3v1024x8m81_1/D
+ pmos_5p0431059130206_3v1024x8m81_0/D pmos_5p0431059130201_3v1024x8m81_0/S pmos_5p0431059130201_3v1024x8m81
Xpmos_5p0431059130209_3v1024x8m81_0 vdd pmos_1p2$$46889004_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ vdd pmos_5p0431059130209_3v1024x8m81_0/S pmos_5p0431059130209_3v1024x8m81
Xpmos_1p2$$46887980_3v1024x8m81_0 vdd vdd pmos_1p2$$46889004_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ pmos_5p0431059130201_3v1024x8m81_0/S pmos_1p2$$46887980_3v1024x8m81
Xpmos_1p2$$46273580_3v1024x8m81_0 pmos_5p0431059130206_3v1024x8m81_0/D men pmos_5p0431059130206_3v1024x8m81_0/D
+ men pmos_1p2$$46273580_3v1024x8m81_0/pmos_5p0431059130203_3v1024x8m81_0/D pmos_5p0431059130206_3v1024x8m81_0/D
+ pmos_1p2$$46273580_3v1024x8m81
Xpmos_5p0431059130206_3v1024x8m81_0 pmos_5p0431059130206_3v1024x8m81_0/D datain pmos_5p0431059130206_3v1024x8m81_0/S
+ pmos_5p0431059130206_3v1024x8m81_0/D nmos_5p04310591302011_3v1024x8m81_1/S pmos_5p0431059130206_3v1024x8m81_0/S
+ pmos_5p0431059130206_3v1024x8m81
Xpmos_1p2$$46273580_3v1024x8m81_1 pmos_5p0431059130206_3v1024x8m81_0/D pmos_5p0431059130201_3v1024x8m81_0/S
+ pmos_5p0431059130206_3v1024x8m81_0/D pmos_5p0431059130201_3v1024x8m81_0/S nmos_5p04310591302011_3v1024x8m81_1/S_uq0
+ pmos_5p0431059130206_3v1024x8m81_0/D pmos_1p2$$46273580_3v1024x8m81
Xnmos_5p04310591302011_3v1024x8m81_0 VSUBS datain pmos_5p0431059130206_3v1024x8m81_0/S
+ nmos_5p04310591302011_3v1024x8m81_1/S pmos_5p0431059130206_3v1024x8m81_0/S VSUBS
+ nmos_5p04310591302011_3v1024x8m81
Xnmos_5p04310591302011_3v1024x8m81_1 nmos_5p04310591302011_3v1024x8m81_1/D pmos_1p2$$46273580_3v1024x8m81_0/pmos_5p0431059130203_3v1024x8m81_0/D
+ men nmos_5p04310591302011_3v1024x8m81_1/S_uq0 nmos_5p04310591302011_3v1024x8m81_1/S
+ VSUBS nmos_5p04310591302011_3v1024x8m81
Xnmos_1p2$$46563372_3v1024x8m81_0 VSUBS nmos_5p04310591302011_3v1024x8m81_1/S_uq0
+ pmos_5p0431059130201_3v1024x8m81_0/S VSUBS nmos_1p2$$46563372_3v1024x8m81
Xnmos_1p2$$46563372_3v1024x8m81_1 VSUBS pmos_1p2$$46273580_3v1024x8m81_0/pmos_5p0431059130203_3v1024x8m81_0/D
+ men VSUBS nmos_1p2$$46563372_3v1024x8m81
Xnmos_5p04310591302010_3v1024x8m81_0 VSUBS nmos_5p04310591302011_3v1024x8m81_1/D pmos_5p0431059130201_3v1024x8m81_0/S
+ VSUBS nmos_5p04310591302010_3v1024x8m81
Xnmos_1p2$$46883884_3v1024x8m81_0 pmos_5p0431059130209_3v1024x8m81_0/S db wep VSUBS
+ nmos_1p2$$46883884_3v1024x8m81
Xnmos_1p2$$46883884_3v1024x8m81_1 VSUBS pmos_5p0431059130209_3v1024x8m81_0/S pmos_1p2$$46889004_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ VSUBS nmos_1p2$$46883884_3v1024x8m81
Xnmos_1p2$$46883884_3v1024x8m81_2 pmos_1p2$$46889004_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ d wep VSUBS nmos_1p2$$46883884_3v1024x8m81
X0 vdd wep a_507_5030# vdd pfet_03v3 ad=0.38572p pd=2.5u as=0.1859p ps=1.23u w=0.695u l=0.28u
X1 a_507_5030# wep vdd vdd pfet_03v3 ad=0.1859p pd=1.23u as=0.38572p ps=2.5u w=0.695u l=0.28u
X2 a_507_5030# wep vss VSUBS nfet_03v3 ad=0.28355p pd=2.13u as=0.3103p ps=2.23u w=0.535u l=0.28u
.ends

.subckt nmos_5p04310591302012_3v1024x8m81 a_n83_n44# D_uq0 D a_77_n44# S_uq1 S_uq0
+ S a_237_n44# a_397_n44# VSUBS
X0 S a_77_n44# D VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.2743p ps=1.575u w=1.055u l=0.28u
X1 S_uq0 a_397_n44# D_uq0 VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D_uq0 a_237_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.2743p ps=1.575u w=1.055u l=0.28u
X3 D a_n83_n44# S_uq1 VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
.ends

.subckt nmos_5p04310591302036_3v1024x8m81 D_uq1 D_uq0 a_530_n44# D a_n112_n44# a_209_n44#
+ a_369_n44# a_48_n44# S_uq1 S_uq0 S VSUBS
X0 D_uq1 a_n112_n44# S_uq1 VSUBS nfet_03v3 ad=0.1378p pd=1.05u as=0.2332p ps=1.94u w=0.53u l=0.28u
X1 S_uq0 a_369_n44# D VSUBS nfet_03v3 ad=0.13913p pd=1.055u as=0.1378p ps=1.05u w=0.53u l=0.28u
X2 D a_209_n44# S VSUBS nfet_03v3 ad=0.1378p pd=1.05u as=0.13913p ps=1.055u w=0.53u l=0.28u
X3 D_uq0 a_530_n44# S_uq0 VSUBS nfet_03v3 ad=0.2332p pd=1.94u as=0.13913p ps=1.055u w=0.53u l=0.28u
X4 S a_48_n44# D_uq1 VSUBS nfet_03v3 ad=0.13913p pd=1.055u as=0.1378p ps=1.05u w=0.53u l=0.28u
.ends

.subckt nmos_1p2$$45101100_3v1024x8m81 nmos_5p04310591302036_3v1024x8m81_0/S a_195_n34#
+ a_35_n34# a_516_n34# nmos_5p04310591302036_3v1024x8m81_0/D nmos_5p04310591302036_3v1024x8m81_0/S_uq1
+ nmos_5p04310591302036_3v1024x8m81_0/S_uq0 a_n125_n34# a_356_n34# nmos_5p04310591302036_3v1024x8m81_0/D_uq1
+ VSUBS nmos_5p04310591302036_3v1024x8m81_0/D_uq0
Xnmos_5p04310591302036_3v1024x8m81_0 nmos_5p04310591302036_3v1024x8m81_0/D_uq1 nmos_5p04310591302036_3v1024x8m81_0/D_uq0
+ a_516_n34# nmos_5p04310591302036_3v1024x8m81_0/D a_n125_n34# a_195_n34# a_356_n34#
+ a_35_n34# nmos_5p04310591302036_3v1024x8m81_0/S_uq1 nmos_5p04310591302036_3v1024x8m81_0/S_uq0
+ nmos_5p04310591302036_3v1024x8m81_0/S VSUBS nmos_5p04310591302036_3v1024x8m81
.ends

.subckt pmos_5p04310591302027_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.28u
.ends

.subckt nmos_5p04310591302033_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1576p pd=1.64u as=0.1576p ps=1.64u w=0.28u l=0.28u
.ends

.subckt pmos_5p04310591302024_3v1024x8m81 w_n286_n86# D_uq1 D_uq0 a_530_n44# D a_n112_n44#
+ a_209_n44# a_369_n44# a_48_n44# S_uq1 S_uq0 S
X0 D_uq1 a_n112_n44# S_uq1 w_n286_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X1 S_uq0 a_369_n44# D w_n286_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D a_209_n44# S w_n286_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.27692p ps=1.58u w=1.055u l=0.28u
X3 D_uq0 a_530_n44# S_uq0 w_n286_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.27692p ps=1.58u w=1.055u l=0.28u
X4 S a_48_n44# D_uq1 w_n286_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46282796_3v1024x8m81 a_n126_n34# pmos_5p04310591302024_3v1024x8m81_0/S_uq1
+ pmos_5p04310591302024_3v1024x8m81_0/S pmos_5p04310591302024_3v1024x8m81_0/S_uq0
+ a_195_n34# pmos_5p04310591302024_3v1024x8m81_0/D_uq1 a_516_n34# pmos_5p04310591302024_3v1024x8m81_0/D_uq0
+ w_163_n66# pmos_5p04310591302024_3v1024x8m81_0/D a_355_n34# a_34_n34#
Xpmos_5p04310591302024_3v1024x8m81_0 w_163_n66# pmos_5p04310591302024_3v1024x8m81_0/D_uq1
+ pmos_5p04310591302024_3v1024x8m81_0/D_uq0 a_516_n34# pmos_5p04310591302024_3v1024x8m81_0/D
+ a_n126_n34# a_195_n34# a_355_n34# a_34_n34# pmos_5p04310591302024_3v1024x8m81_0/S_uq1
+ pmos_5p04310591302024_3v1024x8m81_0/S_uq0 pmos_5p04310591302024_3v1024x8m81_0/S
+ pmos_5p04310591302024_3v1024x8m81
.ends

.subckt pmos_5p04310591302035_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.2067p pd=1.315u as=0.3498p ps=2.47u w=0.795u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.3498p pd=2.47u as=0.2067p ps=1.315u w=0.795u l=0.28u
.ends

.subckt pmos_1p2$$46284844_3v1024x8m81 w_n133_n66# pmos_5p04310591302035_3v1024x8m81_0/S_uq0
+ pmos_5p04310591302035_3v1024x8m81_0/S a_118_n34# a_n42_n34# pmos_5p04310591302035_3v1024x8m81_0/D
Xpmos_5p04310591302035_3v1024x8m81_0 pmos_5p04310591302035_3v1024x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302035_3v1024x8m81_0/S_uq0 pmos_5p04310591302035_3v1024x8m81_0/S
+ pmos_5p04310591302035_3v1024x8m81
.ends

.subckt nmos_5p04310591302023_3v1024x8m81 D a_n32_n44# a_136_n44# S_uq0 S VSUBS
X0 D a_n32_n44# S VSUBS nfet_03v3 ad=92.8f pd=0.92u as=0.1576p ps=1.64u w=0.28u l=0.28u
X1 S_uq0 a_136_n44# D VSUBS nfet_03v3 ad=0.159p pd=1.65u as=92.8f ps=0.92u w=0.28u l=0.28u
.ends

.subckt nmos_5p04310591302029_3v1024x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.54067p pd=3.32u as=0.3159p ps=1.735u w=1.215u l=0.28u
.ends

.subckt nmos_1p2$$45100076_3v1024x8m81 nmos_5p04310591302029_3v1024x8m81_0/D nmos_5p04310591302029_3v1024x8m81_0/S_uq0
+ a_118_n34# a_n41_n34# nmos_5p04310591302029_3v1024x8m81_0/S VSUBS
Xnmos_5p04310591302029_3v1024x8m81_0 nmos_5p04310591302029_3v1024x8m81_0/D a_n41_n34#
+ a_118_n34# nmos_5p04310591302029_3v1024x8m81_0/S_uq0 nmos_5p04310591302029_3v1024x8m81_0/S
+ VSUBS nmos_5p04310591302029_3v1024x8m81
.ends

.subckt nmos_5p04310591302026_3v1024x8m81 D_uq2 D_uq1 D_uq0 a_154_n44# D a_n168_n44#
+ a_476_n44# a_798_n44# a_314_n44# S_uq2 S_uq1 a_n8_n44# S_uq0 S a_636_n44# VSUBS
X0 S_uq0 a_636_n44# D VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
X1 S a_314_n44# D_uq1 VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D_uq2 a_n168_n44# S_uq2 VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X3 S_uq1 a_n8_n44# D_uq2 VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
X4 D_uq0 a_798_n44# S_uq0 VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.27957p ps=1.585u w=1.055u l=0.28u
X5 D a_476_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.27957p ps=1.585u w=1.055u l=0.28u
X6 D_uq1 a_154_n44# S_uq1 VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.27957p ps=1.585u w=1.055u l=0.28u
.ends

.subckt nmos_1p2$$45102124_3v1024x8m81 nmos_5p04310591302026_3v1024x8m81_0/S_uq2 nmos_5p04310591302026_3v1024x8m81_0/S_uq1
+ nmos_5p04310591302026_3v1024x8m81_0/S_uq0 a_140_n34# a_462_n34# nmos_5p04310591302026_3v1024x8m81_0/D_uq2
+ nmos_5p04310591302026_3v1024x8m81_0/S nmos_5p04310591302026_3v1024x8m81_0/D_uq1
+ nmos_5p04310591302026_3v1024x8m81_0/D_uq0 a_n181_n34# a_784_n34# a_300_n34# nmos_5p04310591302026_3v1024x8m81_0/D
+ a_622_n34# a_n22_n34# VSUBS
Xnmos_5p04310591302026_3v1024x8m81_0 nmos_5p04310591302026_3v1024x8m81_0/D_uq2 nmos_5p04310591302026_3v1024x8m81_0/D_uq1
+ nmos_5p04310591302026_3v1024x8m81_0/D_uq0 a_140_n34# nmos_5p04310591302026_3v1024x8m81_0/D
+ a_n181_n34# a_462_n34# a_784_n34# a_300_n34# nmos_5p04310591302026_3v1024x8m81_0/S_uq2
+ nmos_5p04310591302026_3v1024x8m81_0/S_uq1 a_n22_n34# nmos_5p04310591302026_3v1024x8m81_0/S_uq0
+ nmos_5p04310591302026_3v1024x8m81_0/S a_622_n34# VSUBS nmos_5p04310591302026_3v1024x8m81
.ends

.subckt pmos_5p04310591302013_3v1024x8m81 D_uq0 D a_265_n44# S_uq0 S a_n56_n44# a_104_n44#
+ w_n230_n86#
X0 D_uq0 a_265_n44# S_uq0 w_n230_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.27692p ps=1.58u w=1.055u l=0.28u
X1 D a_n56_n44# S w_n230_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X2 S_uq0 a_104_n44# D w_n230_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46286892_3v1024x8m81 w_n133_n66# pmos_5p04310591302013_3v1024x8m81_0/D
+ pmos_5p04310591302013_3v1024x8m81_0/D_uq0 a_251_n34# a_n70_n34# pmos_5p04310591302013_3v1024x8m81_0/S
+ pmos_5p04310591302013_3v1024x8m81_0/S_uq0 a_90_n34#
Xpmos_5p04310591302013_3v1024x8m81_0 pmos_5p04310591302013_3v1024x8m81_0/D_uq0 pmos_5p04310591302013_3v1024x8m81_0/D
+ a_251_n34# pmos_5p04310591302013_3v1024x8m81_0/S_uq0 pmos_5p04310591302013_3v1024x8m81_0/S
+ a_n70_n34# a_90_n34# w_n133_n66# pmos_5p04310591302013_3v1024x8m81
.ends

.subckt pmos_5p04310591302038_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.2464p pd=2u as=0.2464p ps=2u w=0.56u l=0.28u
.ends

.subckt nmos_5p04310591302032_3v1024x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.1378p pd=1.05u as=0.2332p ps=1.94u w=0.53u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.23585p pd=1.95u as=0.1378p ps=1.05u w=0.53u l=0.28u
.ends

.subckt nmos_5p04310591302028_3v1024x8m81 D_uq1 D_uq0 D a_64_n44# a_226_n44# a_386_n44#
+ a_548_n44# S_uq1 S_uq0 S a_n96_n44# VSUBS
X0 D_uq0 a_548_n44# S_uq0 VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.27957p ps=1.585u w=1.055u l=0.28u
X1 S_uq0 a_386_n44# D VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D a_226_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.27957p ps=1.585u w=1.055u l=0.28u
X3 D_uq1 a_n96_n44# S_uq1 VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X4 S a_64_n44# D_uq1 VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_5p04310591302014_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.4642p ps=2.99u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46285868_3v1024x8m81 w_n133_n66# pmos_5p04310591302014_3v1024x8m81_0/S
+ a_n14_n34# pmos_5p04310591302014_3v1024x8m81_0/D
Xpmos_5p04310591302014_3v1024x8m81_0 pmos_5p04310591302014_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302014_3v1024x8m81_0/S pmos_5p04310591302014_3v1024x8m81
.ends

.subckt pmos_5p04310591302031_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.4134p pd=2.11u as=0.6996p ps=4.06u w=1.59u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.6996p pd=4.06u as=0.4134p ps=2.11u w=1.59u l=0.28u
.ends

.subckt pmos_1p2$$46287916_3v1024x8m81 w_n133_n66# a_n42_n34# pmos_5p04310591302031_3v1024x8m81_0/S_uq0
+ pmos_5p04310591302031_3v1024x8m81_0/S a_118_n34# pmos_5p04310591302031_3v1024x8m81_0/D
Xpmos_5p04310591302031_3v1024x8m81_0 pmos_5p04310591302031_3v1024x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302031_3v1024x8m81_0/S_uq0 pmos_5p04310591302031_3v1024x8m81_0/S
+ pmos_5p04310591302031_3v1024x8m81
.ends

.subckt nmos_5p04310591302034_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.2948p pd=2.22u as=0.2948p ps=2.22u w=0.67u l=0.28u
.ends

.subckt pmos_5p04310591302030_3v1024x8m81 D_uq2 a_871_n45# D_uq1 D_uq0 D a_n252_n45#
+ a_550_n45# a_229_n45# w_n426_n86# S_uq4 S_uq2 S_uq3 S_uq1 S_uq0 a_390_n45# S a_n92_n45#
+ a_1032_n45# a_1192_n45# D_uq3 a_711_n45# a_69_n45#
X0 D_uq1 a_390_n45# S_uq2 w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.33205p ps=1.79u w=1.265u l=0.28u
X1 D_uq3 a_n252_n45# S_uq4 w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.5566p ps=3.41u w=1.265u l=0.28u
X2 D_uq2 a_69_n45# S_uq3 w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.33205p ps=1.79u w=1.265u l=0.28u
X3 S_uq2 a_229_n45# D_uq2 w_n426_n86# pfet_03v3 ad=0.33205p pd=1.79u as=0.3289p ps=1.785u w=1.265u l=0.28u
X4 S_uq1 a_550_n45# D_uq1 w_n426_n86# pfet_03v3 ad=0.33205p pd=1.79u as=0.3289p ps=1.785u w=1.265u l=0.28u
X5 S_uq0 a_1192_n45# D_uq0 w_n426_n86# pfet_03v3 ad=0.5566p pd=3.41u as=0.3289p ps=1.785u w=1.265u l=0.28u
X6 D_uq0 a_1032_n45# S w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.33205p ps=1.79u w=1.265u l=0.28u
X7 S_uq3 a_n92_n45# D_uq3 w_n426_n86# pfet_03v3 ad=0.33205p pd=1.79u as=0.3289p ps=1.785u w=1.265u l=0.28u
X8 S a_871_n45# D w_n426_n86# pfet_03v3 ad=0.33205p pd=1.79u as=0.3289p ps=1.785u w=1.265u l=0.28u
X9 D a_711_n45# S_uq1 w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.33205p ps=1.79u w=1.265u l=0.28u
.ends

.subckt pmos_1p2$$45095980_3v1024x8m81 a_697_n34# a_n106_n34# pmos_5p04310591302030_3v1024x8m81_0/S_uq4
+ a_n266_n34# pmos_5p04310591302030_3v1024x8m81_0/S_uq3 a_376_n34# pmos_5p04310591302030_3v1024x8m81_0/S_uq2
+ pmos_5p04310591302030_3v1024x8m81_0/S_uq1 pmos_5p04310591302030_3v1024x8m81_0/S_uq0
+ a_1018_n34# a_1178_n34# pmos_5p04310591302030_3v1024x8m81_0/S a_55_n34# a_857_n34#
+ pmos_5p04310591302030_3v1024x8m81_0/D_uq3 pmos_5p04310591302030_3v1024x8m81_0/D_uq1
+ pmos_5p04310591302030_3v1024x8m81_0/D_uq2 pmos_5p04310591302030_3v1024x8m81_0/D_uq0
+ a_536_n34# w_987_n66# pmos_5p04310591302030_3v1024x8m81_0/D a_215_n34#
Xpmos_5p04310591302030_3v1024x8m81_0 pmos_5p04310591302030_3v1024x8m81_0/D_uq2 a_857_n34#
+ pmos_5p04310591302030_3v1024x8m81_0/D_uq1 pmos_5p04310591302030_3v1024x8m81_0/D_uq0
+ pmos_5p04310591302030_3v1024x8m81_0/D a_n266_n34# a_536_n34# a_215_n34# w_987_n66#
+ pmos_5p04310591302030_3v1024x8m81_0/S_uq4 pmos_5p04310591302030_3v1024x8m81_0/S_uq2
+ pmos_5p04310591302030_3v1024x8m81_0/S_uq3 pmos_5p04310591302030_3v1024x8m81_0/S_uq1
+ pmos_5p04310591302030_3v1024x8m81_0/S_uq0 a_376_n34# pmos_5p04310591302030_3v1024x8m81_0/S
+ a_n106_n34# a_1018_n34# a_1178_n34# pmos_5p04310591302030_3v1024x8m81_0/D_uq3 a_697_n34#
+ a_55_n34# pmos_5p04310591302030_3v1024x8m81
.ends

.subckt pmos_5p04310591302025_3v1024x8m81 D_uq0 D a_265_n44# S_uq0 S a_n56_n44# a_104_n44#
+ w_n230_n85#
X0 D_uq0 a_265_n44# S_uq0 w_n230_n85# pfet_03v3 ad=0.9306p pd=5.11u as=0.55518p ps=2.64u w=2.115u l=0.28u
X1 D a_n56_n44# S w_n230_n85# pfet_03v3 ad=0.5499p pd=2.635u as=0.9306p ps=5.11u w=2.115u l=0.28u
X2 S_uq0 a_104_n44# D w_n230_n85# pfet_03v3 ad=0.55518p pd=2.64u as=0.5499p ps=2.635u w=2.115u l=0.28u
.ends

.subckt pmos_1p2$$46281772_3v1024x8m81 pmos_5p04310591302025_3v1024x8m81_0/D_uq0 pmos_5p04310591302025_3v1024x8m81_0/D
+ a_251_n34# a_n70_n34# w_n133_n66# a_90_n34# pmos_5p04310591302025_3v1024x8m81_0/S_uq0
+ pmos_5p04310591302025_3v1024x8m81_0/S
Xpmos_5p04310591302025_3v1024x8m81_0 pmos_5p04310591302025_3v1024x8m81_0/D_uq0 pmos_5p04310591302025_3v1024x8m81_0/D
+ a_251_n34# pmos_5p04310591302025_3v1024x8m81_0/S_uq0 pmos_5p04310591302025_3v1024x8m81_0/S
+ a_n70_n34# a_90_n34# w_n133_n66# pmos_5p04310591302025_3v1024x8m81
.ends

.subckt nmos_5p04310591302037_3v1024x8m81 a_20_n44# D a_181_n44# a_502_n44# S_uq2
+ a_662_n44# a_n140_n44# S_uq0 a_341_n44# VSUBS
X0 S a_341_n44# D VSUBS nfet_03v3 ad=0.34912p pd=1.855u as=0.3458p ps=1.85u w=1.33u l=0.28u
X1 S_uq0 a_662_n44# D_uq0 VSUBS nfet_03v3 ad=0.5852p pd=3.54u as=0.3458p ps=1.85u w=1.33u l=0.28u
X2 D_uq0 a_502_n44# S VSUBS nfet_03v3 ad=0.3458p pd=1.85u as=0.34912p ps=1.855u w=1.33u l=0.28u
X3 S_uq1 a_20_n44# D_uq1 VSUBS nfet_03v3 ad=0.34912p pd=1.855u as=0.3458p ps=1.85u w=1.33u l=0.28u
X4 D a_181_n44# S_uq1 VSUBS nfet_03v3 ad=0.3458p pd=1.85u as=0.34912p ps=1.855u w=1.33u l=0.28u
X5 D_uq1 a_n140_n44# S_uq2 VSUBS nfet_03v3 ad=0.3458p pd=1.85u as=0.5852p ps=3.54u w=1.33u l=0.28u
.ends

.subckt nmos_1p2$$45103148_3v1024x8m81 a_327_n34# a_n153_n34# nmos_5p04310591302037_3v1024x8m81_0/D
+ nmos_5p04310591302037_3v1024x8m81_0/S_uq2 nmos_5p04310591302037_3v1024x8m81_0/S_uq0
+ a_488_n34# a_167_n34# a_6_n34# a_648_n34# VSUBS
Xnmos_5p04310591302037_3v1024x8m81_0 a_6_n34# nmos_5p04310591302037_3v1024x8m81_0/D
+ a_167_n34# a_488_n34# nmos_5p04310591302037_3v1024x8m81_0/S_uq2 a_648_n34# a_n153_n34#
+ nmos_5p04310591302037_3v1024x8m81_0/S_uq0 a_327_n34# VSUBS nmos_5p04310591302037_3v1024x8m81
.ends

.subckt pmos_5p04310591302022_3v1024x8m81 D_uq2 D_uq1 D_uq0 D a_n252_n44# a_550_n44#
+ a_229_n44# w_n426_n86# S_uq4 S_uq2 S_uq3 S_uq1 a_390_n44# S_uq0 S a_n92_n44# a_1032_n44#
+ a_1192_n44# a_711_n44# a_69_n44# D_uq3 a_871_n44#
X0 D_uq1 a_390_n44# S_uq2 w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.50005p ps=2.43u w=1.905u l=0.28u
X1 D_uq3 a_n252_n44# S_uq4 w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.8382p ps=4.69u w=1.905u l=0.28u
X2 D_uq2 a_69_n44# S_uq3 w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.50005p ps=2.43u w=1.905u l=0.28u
X3 S_uq2 a_229_n44# D_uq2 w_n426_n86# pfet_03v3 ad=0.50005p pd=2.43u as=0.4953p ps=2.425u w=1.905u l=0.28u
X4 S_uq1 a_550_n44# D_uq1 w_n426_n86# pfet_03v3 ad=0.50005p pd=2.43u as=0.4953p ps=2.425u w=1.905u l=0.28u
X5 S_uq0 a_1192_n44# D_uq0 w_n426_n86# pfet_03v3 ad=0.8382p pd=4.69u as=0.4953p ps=2.425u w=1.905u l=0.28u
X6 D_uq0 a_1032_n44# S w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.50005p ps=2.43u w=1.905u l=0.28u
X7 S_uq3 a_n92_n44# D_uq3 w_n426_n86# pfet_03v3 ad=0.50005p pd=2.43u as=0.4953p ps=2.425u w=1.905u l=0.28u
X8 S a_871_n44# D w_n426_n86# pfet_03v3 ad=0.50005p pd=2.43u as=0.4953p ps=2.425u w=1.905u l=0.28u
X9 D a_711_n44# S_uq1 w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.50005p ps=2.43u w=1.905u l=0.28u
.ends

.subckt pmos_1p2$$46283820_3v1024x8m81 a_536_n34# a_215_n34# a_697_n34# pmos_5p04310591302022_3v1024x8m81_0/S_uq3
+ pmos_5p04310591302022_3v1024x8m81_0/S_uq4 pmos_5p04310591302022_3v1024x8m81_0/S_uq2
+ a_n106_n34# pmos_5p04310591302022_3v1024x8m81_0/S_uq1 a_n266_n34# pmos_5p04310591302022_3v1024x8m81_0/S_uq0
+ pmos_5p04310591302022_3v1024x8m81_0/S a_376_n34# w_984_n66# a_1018_n34# a_1178_n34#
+ a_55_n34# pmos_5p04310591302022_3v1024x8m81_0/D_uq3 pmos_5p04310591302022_3v1024x8m81_0/D_uq2
+ pmos_5p04310591302022_3v1024x8m81_0/D_uq1 a_857_n34# pmos_5p04310591302022_3v1024x8m81_0/D_uq0
+ pmos_5p04310591302022_3v1024x8m81_0/D
Xpmos_5p04310591302022_3v1024x8m81_0 pmos_5p04310591302022_3v1024x8m81_0/D_uq2 pmos_5p04310591302022_3v1024x8m81_0/D_uq1
+ pmos_5p04310591302022_3v1024x8m81_0/D_uq0 pmos_5p04310591302022_3v1024x8m81_0/D
+ a_n266_n34# a_536_n34# a_215_n34# w_984_n66# pmos_5p04310591302022_3v1024x8m81_0/S_uq4
+ pmos_5p04310591302022_3v1024x8m81_0/S_uq2 pmos_5p04310591302022_3v1024x8m81_0/S_uq3
+ pmos_5p04310591302022_3v1024x8m81_0/S_uq1 a_376_n34# pmos_5p04310591302022_3v1024x8m81_0/S_uq0
+ pmos_5p04310591302022_3v1024x8m81_0/S a_n106_n34# a_1018_n34# a_1178_n34# a_697_n34#
+ a_55_n34# pmos_5p04310591302022_3v1024x8m81_0/D_uq3 a_857_n34# pmos_5p04310591302022_3v1024x8m81
.ends

.subckt sacntl_2_3v1024x8m81 pcb se pmos_5p04310591302027_3v1024x8m81_1/S_uq0 men
+ pmos_5p04310591302027_3v1024x8m81_2/S_uq0 vdd vdd_uq0 vss
Xnmos_5p04310591302012_3v1024x8m81_0 nmos_5p04310591302028_3v1024x8m81_1/S se se nmos_5p04310591302028_3v1024x8m81_1/S
+ vss vss vss nmos_5p04310591302028_3v1024x8m81_1/S nmos_5p04310591302028_3v1024x8m81_1/S
+ vss nmos_5p04310591302012_3v1024x8m81
Xnmos_1p2$$45101100_3v1024x8m81_0 vss men men men pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D
+ vss vss men men pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D
+ vss pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D nmos_1p2$$45101100_3v1024x8m81
Xpmos_5p04310591302027_3v1024x8m81_0 vdd_uq0 pmos_5p04310591302027_3v1024x8m81_2/S_uq0
+ pmos_5p04310591302027_3v1024x8m81_0/S vdd_uq0 pmos_5p04310591302027_3v1024x8m81_0/S_uq0
+ pmos_5p04310591302027_3v1024x8m81_0/S pmos_5p04310591302027_3v1024x8m81
Xnmos_5p04310591302033_3v1024x8m81_0 vss pmos_5p04310591302027_3v1024x8m81_0/S_uq0
+ pmos_5p04310591302038_3v1024x8m81_0/S vss nmos_5p04310591302033_3v1024x8m81
Xpmos_5p04310591302027_3v1024x8m81_1 vdd_uq0 pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D
+ vss vdd_uq0 pmos_5p04310591302027_3v1024x8m81_1/S_uq0 pmos_5p04310591302027_3v1024x8m81_1/S
+ pmos_5p04310591302027_3v1024x8m81
Xpmos_5p04310591302027_3v1024x8m81_2 vdd_uq0 pmos_5p04310591302027_3v1024x8m81_1/S_uq0
+ pmos_5p04310591302027_3v1024x8m81_2/S vdd_uq0 pmos_5p04310591302027_3v1024x8m81_2/S_uq0
+ pmos_5p04310591302027_3v1024x8m81_2/S pmos_5p04310591302027_3v1024x8m81
Xpmos_1p2$$46282796_3v1024x8m81_0 men vdd_uq0 vdd_uq0 vdd_uq0 men pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D
+ men pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D vdd_uq0
+ pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D men men pmos_1p2$$46282796_3v1024x8m81
Xpmos_1p2$$46284844_3v1024x8m81_0 vdd_uq0 vdd_uq0 vdd_uq0 pmos_5p04310591302027_3v1024x8m81_1/S
+ pmos_5p04310591302027_3v1024x8m81_1/S nmos_5p04310591302034_3v1024x8m81_0/D pmos_1p2$$46284844_3v1024x8m81
Xnmos_5p04310591302023_3v1024x8m81_0 vss pmos_5p04310591302027_3v1024x8m81_2/S_uq0
+ pmos_5p04310591302027_3v1024x8m81_0/S pmos_5p04310591302027_3v1024x8m81_0/S_uq0
+ pmos_5p04310591302027_3v1024x8m81_0/S vss nmos_5p04310591302023_3v1024x8m81
Xnmos_1p2$$45100076_3v1024x8m81_0 pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S
+ vss pmos_1p2$$46281772_3v1024x8m81_1/pmos_5p04310591302025_3v1024x8m81_0/S pmos_1p2$$46281772_3v1024x8m81_1/pmos_5p04310591302025_3v1024x8m81_0/S
+ vss vss nmos_1p2$$45100076_3v1024x8m81
Xnmos_5p04310591302023_3v1024x8m81_1 vss pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D
+ vss pmos_5p04310591302027_3v1024x8m81_1/S_uq0 pmos_5p04310591302027_3v1024x8m81_1/S
+ vss nmos_5p04310591302023_3v1024x8m81
Xnmos_5p04310591302023_3v1024x8m81_2 vss pmos_5p04310591302027_3v1024x8m81_1/S_uq0
+ pmos_5p04310591302027_3v1024x8m81_2/S pmos_5p04310591302027_3v1024x8m81_2/S_uq0
+ pmos_5p04310591302027_3v1024x8m81_2/S vss nmos_5p04310591302023_3v1024x8m81
Xnmos_1p2$$45102124_3v1024x8m81_0 vss vss vss pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S
+ pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S pcb vss pcb
+ pcb pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S
+ pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S pcb pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S
+ pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S vss nmos_1p2$$45102124_3v1024x8m81
Xpmos_1p2$$46286892_3v1024x8m81_0 vdd nmos_5p04310591302028_3v1024x8m81_1/S nmos_5p04310591302028_3v1024x8m81_1/S
+ nmos_5p04310591302032_3v1024x8m81_0/D nmos_5p04310591302032_3v1024x8m81_0/D vdd
+ vdd nmos_5p04310591302032_3v1024x8m81_0/D pmos_1p2$$46286892_3v1024x8m81
Xpmos_5p04310591302038_3v1024x8m81_0 vdd_uq0 pmos_5p04310591302027_3v1024x8m81_0/S_uq0
+ vdd_uq0 pmos_5p04310591302038_3v1024x8m81_0/S pmos_5p04310591302038_3v1024x8m81
Xnmos_5p04310591302032_3v1024x8m81_0 nmos_5p04310591302032_3v1024x8m81_0/D nmos_5p04310591302034_3v1024x8m81_0/D
+ nmos_5p04310591302034_3v1024x8m81_0/D vss vss vss nmos_5p04310591302032_3v1024x8m81
Xnmos_5p04310591302028_3v1024x8m81_0 nmos_5p04310591302028_3v1024x8m81_1/D nmos_5p04310591302028_3v1024x8m81_1/D
+ nmos_5p04310591302028_3v1024x8m81_1/D nmos_5p04310591302032_3v1024x8m81_0/D nmos_5p04310591302032_3v1024x8m81_0/D
+ nmos_5p04310591302032_3v1024x8m81_0/D nmos_5p04310591302032_3v1024x8m81_0/D vss
+ vss vss nmos_5p04310591302032_3v1024x8m81_0/D vss nmos_5p04310591302028_3v1024x8m81
Xnmos_5p04310591302028_3v1024x8m81_1 nmos_5p04310591302028_3v1024x8m81_1/D nmos_5p04310591302028_3v1024x8m81_1/D
+ nmos_5p04310591302028_3v1024x8m81_1/D pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D
+ pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D
+ pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D nmos_5p04310591302028_3v1024x8m81_1/S
+ nmos_5p04310591302028_3v1024x8m81_1/S nmos_5p04310591302028_3v1024x8m81_1/S pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D
+ vss nmos_5p04310591302028_3v1024x8m81
Xpmos_1p2$$46285868_3v1024x8m81_0 vdd nmos_5p04310591302028_3v1024x8m81_1/S pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D
+ vdd pmos_1p2$$46285868_3v1024x8m81
Xpmos_1p2$$46287916_3v1024x8m81_0 vdd nmos_5p04310591302034_3v1024x8m81_0/D vdd vdd
+ nmos_5p04310591302034_3v1024x8m81_0/D nmos_5p04310591302032_3v1024x8m81_0/D pmos_1p2$$46287916_3v1024x8m81
Xnmos_5p04310591302034_3v1024x8m81_0 nmos_5p04310591302034_3v1024x8m81_0/D pmos_5p04310591302027_3v1024x8m81_1/S
+ vss vss nmos_5p04310591302034_3v1024x8m81
Xpmos_1p2$$45095980_3v1024x8m81_0 nmos_5p04310591302028_3v1024x8m81_1/S nmos_5p04310591302028_3v1024x8m81_1/S
+ vdd nmos_5p04310591302028_3v1024x8m81_1/S vdd nmos_5p04310591302028_3v1024x8m81_1/S
+ vdd vdd vdd nmos_5p04310591302028_3v1024x8m81_1/S nmos_5p04310591302028_3v1024x8m81_1/S
+ vdd nmos_5p04310591302028_3v1024x8m81_1/S nmos_5p04310591302028_3v1024x8m81_1/S
+ se se se se nmos_5p04310591302028_3v1024x8m81_1/S vdd se nmos_5p04310591302028_3v1024x8m81_1/S
+ pmos_1p2$$45095980_3v1024x8m81
Xpmos_1p2$$46281772_3v1024x8m81_0 vdd vdd pmos_1p2$$46281772_3v1024x8m81_1/pmos_5p04310591302025_3v1024x8m81_0/S
+ pmos_1p2$$46281772_3v1024x8m81_1/pmos_5p04310591302025_3v1024x8m81_0/S vdd pmos_1p2$$46281772_3v1024x8m81_1/pmos_5p04310591302025_3v1024x8m81_0/S
+ pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S
+ pmos_1p2$$46281772_3v1024x8m81
Xpmos_1p2$$46281772_3v1024x8m81_1 vdd vdd nmos_5p04310591302028_3v1024x8m81_1/S pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D
+ vdd nmos_5p04310591302034_3v1024x8m81_0/D pmos_1p2$$46281772_3v1024x8m81_1/pmos_5p04310591302025_3v1024x8m81_0/S
+ pmos_1p2$$46281772_3v1024x8m81_1/pmos_5p04310591302025_3v1024x8m81_0/S pmos_1p2$$46281772_3v1024x8m81
Xnmos_1p2$$45103148_3v1024x8m81_0 nmos_5p04310591302028_3v1024x8m81_1/S pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D
+ pmos_1p2$$46281772_3v1024x8m81_1/pmos_5p04310591302025_3v1024x8m81_0/S vss vss nmos_5p04310591302034_3v1024x8m81_0/D
+ nmos_5p04310591302028_3v1024x8m81_1/S nmos_5p04310591302034_3v1024x8m81_0/D pmos_1p2$$46282796_3v1024x8m81_0/pmos_5p04310591302024_3v1024x8m81_0/D
+ vss nmos_1p2$$45103148_3v1024x8m81
Xpmos_1p2$$46283820_3v1024x8m81_0 pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S
+ pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S
+ vdd vdd vdd pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S
+ vdd pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S vdd vdd
+ pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S vdd pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S
+ pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S
+ pcb pcb pcb pmos_1p2$$46281772_3v1024x8m81_0/pmos_5p04310591302025_3v1024x8m81_0/S
+ pcb pcb pmos_1p2$$46283820_3v1024x8m81
.ends

.subckt nmos_5p04310591302016_3v1024x8m81 D_uq2 a_124_n45# D_uq1 a_284_n45# D_uq0
+ D a_446_n45# a_768_n45# a_n198_n45# a_n38_n45# S_uq2 S_uq3 S_uq1 S_uq0 a_606_n45#
+ S a_928_n45# VSUBS
X0 S_uq0 a_928_n45# D_uq0 VSUBS nfet_03v3 ad=0.7155p pd=4.08u as=0.4134p ps=2.11u w=1.59u l=0.28u
X1 D_uq2 a_n198_n45# S_uq3 VSUBS nfet_03v3 ad=0.4134p pd=2.11u as=0.70755p ps=4.07u w=1.59u l=0.28u
X2 S_uq2 a_n38_n45# D_uq2 VSUBS nfet_03v3 ad=0.42135p pd=2.12u as=0.4134p ps=2.11u w=1.59u l=0.28u
X3 S a_606_n45# D VSUBS nfet_03v3 ad=0.42135p pd=2.12u as=0.4134p ps=2.11u w=1.59u l=0.28u
X4 D_uq0 a_768_n45# S VSUBS nfet_03v3 ad=0.4134p pd=2.11u as=0.42135p ps=2.12u w=1.59u l=0.28u
X5 D a_446_n45# S_uq1 VSUBS nfet_03v3 ad=0.4134p pd=2.11u as=0.42135p ps=2.12u w=1.59u l=0.28u
X6 S_uq1 a_284_n45# D_uq1 VSUBS nfet_03v3 ad=0.42135p pd=2.12u as=0.4134p ps=2.11u w=1.59u l=0.28u
X7 D_uq1 a_124_n45# S_uq2 VSUBS nfet_03v3 ad=0.4134p pd=2.11u as=0.42135p ps=2.12u w=1.59u l=0.28u
.ends

.subckt nmos_1p2$$46552108_3v1024x8m81 nmos_5p04310591302016_3v1024x8m81_0/a_124_n45#
+ nmos_5p04310591302016_3v1024x8m81_0/a_284_n45# nmos_5p04310591302016_3v1024x8m81_0/a_446_n45#
+ nmos_5p04310591302016_3v1024x8m81_0/D nmos_5p04310591302016_3v1024x8m81_0/a_768_n45#
+ nmos_5p04310591302016_3v1024x8m81_0/a_n198_n45# nmos_5p04310591302016_3v1024x8m81_0/a_n38_n45#
+ nmos_5p04310591302016_3v1024x8m81_0/S_uq3 nmos_5p04310591302016_3v1024x8m81_0/S_uq1
+ nmos_5p04310591302016_3v1024x8m81_0/S_uq2 nmos_5p04310591302016_3v1024x8m81_0/S_uq0
+ nmos_5p04310591302016_3v1024x8m81_0/a_606_n45# nmos_5p04310591302016_3v1024x8m81_0/S
+ nmos_5p04310591302016_3v1024x8m81_0/a_928_n45# nmos_5p04310591302016_3v1024x8m81_0/D_uq2
+ nmos_5p04310591302016_3v1024x8m81_0/D_uq1 VSUBS nmos_5p04310591302016_3v1024x8m81_0/D_uq0
Xnmos_5p04310591302016_3v1024x8m81_0 nmos_5p04310591302016_3v1024x8m81_0/D_uq2 nmos_5p04310591302016_3v1024x8m81_0/a_124_n45#
+ nmos_5p04310591302016_3v1024x8m81_0/D_uq1 nmos_5p04310591302016_3v1024x8m81_0/a_284_n45#
+ nmos_5p04310591302016_3v1024x8m81_0/D_uq0 nmos_5p04310591302016_3v1024x8m81_0/D
+ nmos_5p04310591302016_3v1024x8m81_0/a_446_n45# nmos_5p04310591302016_3v1024x8m81_0/a_768_n45#
+ nmos_5p04310591302016_3v1024x8m81_0/a_n198_n45# nmos_5p04310591302016_3v1024x8m81_0/a_n38_n45#
+ nmos_5p04310591302016_3v1024x8m81_0/S_uq2 nmos_5p04310591302016_3v1024x8m81_0/S_uq3
+ nmos_5p04310591302016_3v1024x8m81_0/S_uq1 nmos_5p04310591302016_3v1024x8m81_0/S_uq0
+ nmos_5p04310591302016_3v1024x8m81_0/a_606_n45# nmos_5p04310591302016_3v1024x8m81_0/S
+ nmos_5p04310591302016_3v1024x8m81_0/a_928_n45# VSUBS nmos_5p04310591302016_3v1024x8m81
.ends

.subckt nmos_1p2$$45107244_3v1024x8m81 nmos_5p04310591302012_3v1024x8m81_0/D a_223_n34#
+ a_383_n34# nmos_5p04310591302012_3v1024x8m81_0/S_uq1 nmos_5p04310591302012_3v1024x8m81_0/S_uq0
+ nmos_5p04310591302012_3v1024x8m81_0/S a_n96_n34# nmos_5p04310591302012_3v1024x8m81_0/D_uq0
+ a_63_n34# VSUBS
Xnmos_5p04310591302012_3v1024x8m81_0 a_n96_n34# nmos_5p04310591302012_3v1024x8m81_0/D_uq0
+ nmos_5p04310591302012_3v1024x8m81_0/D a_63_n34# nmos_5p04310591302012_3v1024x8m81_0/S_uq1
+ nmos_5p04310591302012_3v1024x8m81_0/S_uq0 nmos_5p04310591302012_3v1024x8m81_0/S
+ a_223_n34# a_383_n34# VSUBS nmos_5p04310591302012_3v1024x8m81
.ends

.subckt pmos_5p04310591302021_3v1024x8m81 a_76_n44# D_uq0 D a_n84_n44# w_n258_n86#
+ S_uq1 S_uq0 S a_237_n44# a_397_n44#
X0 S_uq0 a_397_n44# D_uq0 w_n258_n86# pfet_03v3 ad=0.1848p pd=1.72u as=0.1092p ps=0.94u w=0.42u l=0.28u
X1 D_uq0 a_237_n44# S w_n258_n86# pfet_03v3 ad=0.1092p pd=0.94u as=0.11025p ps=0.945u w=0.42u l=0.28u
X2 D a_n84_n44# S_uq1 w_n258_n86# pfet_03v3 ad=0.1092p pd=0.94u as=0.1848p ps=1.72u w=0.42u l=0.28u
X3 S a_76_n44# D w_n258_n86# pfet_03v3 ad=0.11025p pd=0.945u as=0.1092p ps=0.94u w=0.42u l=0.28u
.ends

.subckt pmos_1p2$$46896172_3v1024x8m81 w_n133_n66# pmos_5p04310591302021_3v1024x8m81_0/D_uq0
+ pmos_5p04310591302021_3v1024x8m81_0/D pmos_5p04310591302021_3v1024x8m81_0/a_n84_n44#
+ pmos_5p04310591302021_3v1024x8m81_0/S_uq1 pmos_5p04310591302021_3v1024x8m81_0/S_uq0
+ pmos_5p04310591302021_3v1024x8m81_0/S pmos_5p04310591302021_3v1024x8m81_0/a_237_n44#
+ pmos_5p04310591302021_3v1024x8m81_0/a_397_n44# pmos_5p04310591302021_3v1024x8m81_0/a_76_n44#
Xpmos_5p04310591302021_3v1024x8m81_0 pmos_5p04310591302021_3v1024x8m81_0/a_76_n44#
+ pmos_5p04310591302021_3v1024x8m81_0/D_uq0 pmos_5p04310591302021_3v1024x8m81_0/D
+ pmos_5p04310591302021_3v1024x8m81_0/a_n84_n44# w_n133_n66# pmos_5p04310591302021_3v1024x8m81_0/S_uq1
+ pmos_5p04310591302021_3v1024x8m81_0/S_uq0 pmos_5p04310591302021_3v1024x8m81_0/S
+ pmos_5p04310591302021_3v1024x8m81_0/a_237_n44# pmos_5p04310591302021_3v1024x8m81_0/a_397_n44#
+ pmos_5p04310591302021_3v1024x8m81
.ends

.subckt pmos_5p04310591302019_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.1848p pd=1.72u as=0.1848p ps=1.72u w=0.42u l=0.28u
.ends

.subckt pmos_1p2$$46898220_3v1024x8m81 w_n133_n66# pmos_5p04310591302019_3v1024x8m81_0/D
+ a_n14_84# pmos_5p04310591302019_3v1024x8m81_0/S
Xpmos_5p04310591302019_3v1024x8m81_0 pmos_5p04310591302019_3v1024x8m81_0/D a_n14_84#
+ w_n133_n66# pmos_5p04310591302019_3v1024x8m81_0/S pmos_5p04310591302019_3v1024x8m81
.ends

.subckt pmos_5p04310591302018_3v1024x8m81 D_uq1 a_20_n45# D_uq0 D a_181_n45# S_uq2
+ a_502_n45# S_uq1 a_662_n45# a_n140_n45# S_uq0 S a_341_n45# w_n314_n86#
X0 S a_341_n45# D w_n314_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
X1 S_uq0 a_662_n45# D_uq0 w_n314_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D_uq0 a_502_n45# S w_n314_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.27692p ps=1.58u w=1.055u l=0.28u
X3 S_uq1 a_20_n45# D_uq1 w_n314_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
X4 D a_181_n45# S_uq1 w_n314_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.27692p ps=1.58u w=1.055u l=0.28u
X5 D_uq1 a_n140_n45# S_uq2 w_n314_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46549036_3v1024x8m81 a_327_n34# w_n188_n50# pmos_5p04310591302018_3v1024x8m81_0/D
+ pmos_5p04310591302018_3v1024x8m81_0/D_uq0 pmos_5p04310591302018_3v1024x8m81_0/D_uq1
+ a_488_n34# a_n154_n34# a_167_n34# a_6_n34# pmos_5p04310591302018_3v1024x8m81_0/S
+ a_648_n34# pmos_5p04310591302018_3v1024x8m81_0/S_uq2 pmos_5p04310591302018_3v1024x8m81_0/S_uq1
+ pmos_5p04310591302018_3v1024x8m81_0/S_uq0
Xpmos_5p04310591302018_3v1024x8m81_0 pmos_5p04310591302018_3v1024x8m81_0/D_uq1 a_6_n34#
+ pmos_5p04310591302018_3v1024x8m81_0/D_uq0 pmos_5p04310591302018_3v1024x8m81_0/D
+ a_167_n34# pmos_5p04310591302018_3v1024x8m81_0/S_uq2 a_488_n34# pmos_5p04310591302018_3v1024x8m81_0/S_uq1
+ a_648_n34# a_n154_n34# pmos_5p04310591302018_3v1024x8m81_0/S_uq0 pmos_5p04310591302018_3v1024x8m81_0/S
+ a_327_n34# w_n188_n50# pmos_5p04310591302018_3v1024x8m81
.ends

.subckt nmos_5p04310591302017_3v1024x8m81 D_uq2 D_uq1 a_n37_n44# D_uq0 D a_929_n44#
+ a_125_n44# a_285_n44# a_447_n44# a_769_n44# S_uq2 S_uq3 S_uq1 S_uq0 S a_607_n44#
+ a_n197_n44# VSUBS
X0 D_uq0 a_769_n44# S VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.35112p ps=1.855u w=1.325u l=0.28u
X1 D a_447_n44# S_uq1 VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.35112p ps=1.855u w=1.325u l=0.28u
X2 D_uq2 a_n197_n44# S_uq3 VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.583p ps=3.53u w=1.325u l=0.28u
X3 S_uq2 a_n37_n44# D_uq2 VSUBS nfet_03v3 ad=0.35112p pd=1.855u as=0.3445p ps=1.845u w=1.325u l=0.28u
X4 S_uq1 a_285_n44# D_uq1 VSUBS nfet_03v3 ad=0.35112p pd=1.855u as=0.3445p ps=1.845u w=1.325u l=0.28u
X5 D_uq1 a_125_n44# S_uq2 VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.35112p ps=1.855u w=1.325u l=0.28u
X6 S_uq0 a_929_n44# D_uq0 VSUBS nfet_03v3 ad=0.58963p pd=3.54u as=0.3445p ps=1.845u w=1.325u l=0.28u
X7 S a_607_n44# D VSUBS nfet_03v3 ad=0.35112p pd=1.855u as=0.3445p ps=1.845u w=1.325u l=0.28u
.ends

.subckt nmos_1p2$$46550060_3v1024x8m81 nmos_5p04310591302017_3v1024x8m81_0/D a_915_n34#
+ nmos_5p04310591302017_3v1024x8m81_0/S_uq3 nmos_5p04310591302017_3v1024x8m81_0/S_uq2
+ nmos_5p04310591302017_3v1024x8m81_0/S_uq1 nmos_5p04310591302017_3v1024x8m81_0/S_uq0
+ a_111_n34# a_271_n34# a_433_n34# nmos_5p04310591302017_3v1024x8m81_0/S a_593_n34#
+ a_n51_n34# a_755_n34# nmos_5p04310591302017_3v1024x8m81_0/D_uq2 nmos_5p04310591302017_3v1024x8m81_0/D_uq1
+ a_n210_n34# nmos_5p04310591302017_3v1024x8m81_0/D_uq0 VSUBS
Xnmos_5p04310591302017_3v1024x8m81_0 nmos_5p04310591302017_3v1024x8m81_0/D_uq2 nmos_5p04310591302017_3v1024x8m81_0/D_uq1
+ a_n51_n34# nmos_5p04310591302017_3v1024x8m81_0/D_uq0 nmos_5p04310591302017_3v1024x8m81_0/D
+ a_915_n34# a_111_n34# a_271_n34# a_433_n34# a_755_n34# nmos_5p04310591302017_3v1024x8m81_0/S_uq2
+ nmos_5p04310591302017_3v1024x8m81_0/S_uq3 nmos_5p04310591302017_3v1024x8m81_0/S_uq1
+ nmos_5p04310591302017_3v1024x8m81_0/S_uq0 nmos_5p04310591302017_3v1024x8m81_0/S
+ a_593_n34# a_n210_n34# VSUBS nmos_5p04310591302017_3v1024x8m81
.ends

.subckt pmos_5p04310591302020_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46897196_3v1024x8m81 w_n133_n66# a_n42_n34# pmos_5p04310591302020_3v1024x8m81_0/D
+ a_118_n34# pmos_5p04310591302020_3v1024x8m81_0/S_uq0 pmos_5p04310591302020_3v1024x8m81_0/S
Xpmos_5p04310591302020_3v1024x8m81_0 pmos_5p04310591302020_3v1024x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302020_3v1024x8m81_0/S_uq0 pmos_5p04310591302020_3v1024x8m81_0/S
+ pmos_5p04310591302020_3v1024x8m81
.ends

.subckt nmos_1p2$$46551084_3v1024x8m81 nmos_5p04310591302010_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v1024x8m81_0/S VSUBS
Xnmos_5p04310591302010_3v1024x8m81_0 nmos_5p04310591302010_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v1024x8m81_0/S VSUBS nmos_5p04310591302010_3v1024x8m81
.ends

.subckt nmos_5p04310591302015_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.6996p pd=4.06u as=0.6996p ps=4.06u w=1.59u l=0.28u
.ends

.subckt nmos_1p2$$46553132_3v1024x8m81 nmos_5p04310591302015_3v1024x8m81_0/S nmos_5p04310591302015_3v1024x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p04310591302015_3v1024x8m81_0 nmos_5p04310591302015_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p04310591302015_3v1024x8m81_0/S VSUBS nmos_5p04310591302015_3v1024x8m81
.ends

.subckt sa_3v1024x8m81 qp qn wep se pcb db pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D
+ vdd d vss
Xnmos_1p2$$46552108_3v1024x8m81_0 pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D
+ pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S
+ nmos_1p2$$46552108_3v1024x8m81_0/nmos_5p04310591302016_3v1024x8m81_0/D pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D
+ pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D
+ pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D
+ pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D
+ pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S
+ pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S nmos_1p2$$46552108_3v1024x8m81_0/nmos_5p04310591302016_3v1024x8m81_0/D
+ nmos_1p2$$46552108_3v1024x8m81_0/nmos_5p04310591302016_3v1024x8m81_0/D vss nmos_1p2$$46552108_3v1024x8m81_0/nmos_5p04310591302016_3v1024x8m81_0/D
+ nmos_1p2$$46552108_3v1024x8m81
Xnmos_1p2$$45107244_3v1024x8m81_0 vss nmos_1p2$$46551084_3v1024x8m81_0/nmos_5p04310591302010_3v1024x8m81_0/S
+ nmos_1p2$$46551084_3v1024x8m81_0/nmos_5p04310591302010_3v1024x8m81_0/S qn qp qp
+ pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D vss nmos_1p2$$46551084_3v1024x8m81_0/nmos_5p04310591302010_3v1024x8m81_0/S
+ vss nmos_1p2$$45107244_3v1024x8m81
Xpmos_1p2$$46896172_3v1024x8m81_0 pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D
+ pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D
+ pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S
+ pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D
+ pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D
+ pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S pmos_1p2$$46896172_3v1024x8m81
Xpmos_1p2$$46898220_3v1024x8m81_0 pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D
+ pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D
+ pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D pmos_1p2$$46898220_3v1024x8m81
Xpmos_1p2$$46898220_3v1024x8m81_1 pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D
+ pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D
+ pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S pmos_1p2$$46898220_3v1024x8m81
Xpmos_1p2$$46549036_3v1024x8m81_0 nmos_1p2$$46551084_3v1024x8m81_0/nmos_5p04310591302010_3v1024x8m81_0/S
+ vdd qp nmos_1p2$$46551084_3v1024x8m81_0/nmos_5p04310591302010_3v1024x8m81_0/S qn
+ pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D
+ nmos_1p2$$46551084_3v1024x8m81_0/nmos_5p04310591302010_3v1024x8m81_0/S pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D
+ vdd pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S vdd vdd
+ vdd pmos_1p2$$46549036_3v1024x8m81
Xnmos_1p2$$46550060_3v1024x8m81_0 nmos_1p2$$46552108_3v1024x8m81_0/nmos_5p04310591302016_3v1024x8m81_0/D
+ se vss vss vss vss se se se vss se se se nmos_1p2$$46552108_3v1024x8m81_0/nmos_5p04310591302016_3v1024x8m81_0/D
+ nmos_1p2$$46552108_3v1024x8m81_0/nmos_5p04310591302016_3v1024x8m81_0/D se nmos_1p2$$46552108_3v1024x8m81_0/nmos_5p04310591302016_3v1024x8m81_0/D
+ vss nmos_1p2$$46550060_3v1024x8m81
Xpmos_1p2$$46286892_3v1024x8m81_0 pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D
+ d pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D pcb pcb
+ pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D db pcb pmos_1p2$$46286892_3v1024x8m81
Xpmos_1p2$$46897196_3v1024x8m81_0 pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D
+ se pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S se d d
+ pmos_1p2$$46897196_3v1024x8m81
Xpmos_1p2$$46897196_3v1024x8m81_1 pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D
+ se pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D se db
+ db pmos_1p2$$46897196_3v1024x8m81
Xpmos_1p2$$46897196_3v1024x8m81_2 pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D
+ se pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D se db
+ db pmos_1p2$$46897196_3v1024x8m81
Xpmos_1p2$$46285868_3v1024x8m81_0 pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D
+ pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D pcb pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S
+ pmos_1p2$$46285868_3v1024x8m81
Xpmos_1p2$$46897196_3v1024x8m81_3 pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/D
+ se pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S se d d
+ pmos_1p2$$46897196_3v1024x8m81
Xnmos_1p2$$46551084_3v1024x8m81_0 vss pmos_1p2$$46898220_3v1024x8m81_1/pmos_5p04310591302019_3v1024x8m81_0/S
+ nmos_1p2$$46551084_3v1024x8m81_0/nmos_5p04310591302010_3v1024x8m81_0/S vss nmos_1p2$$46551084_3v1024x8m81
Xnmos_1p2$$46553132_3v1024x8m81_0 pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D
+ vss vss vss nmos_1p2$$46553132_3v1024x8m81
Xnmos_1p2$$46553132_3v1024x8m81_1 vss pmos_1p2$$46897196_3v1024x8m81_2/pmos_5p04310591302020_3v1024x8m81_0/D
+ vss vss nmos_1p2$$46553132_3v1024x8m81
.ends

.subckt nmos_5p0431059130200_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.397p pd=7.23u as=1.397p ps=7.23u w=3.175u l=0.28u
.ends

.subckt nmos_1p2$$47119404_3v1024x8m81 nmos_5p0431059130200_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p0431059130200_3v1024x8m81_0/S VSUBS
Xnmos_5p0431059130200_3v1024x8m81_0 nmos_5p0431059130200_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p0431059130200_3v1024x8m81_0/S VSUBS nmos_5p0431059130200_3v1024x8m81
.ends

.subckt nmos_5p0431059130202_3v1024x8m81 D a_n32_n44# a_136_n44# S_uq0 S VSUBS
X0 D a_n32_n44# S VSUBS nfet_03v3 ad=91.3f pd=0.92u as=0.1561p ps=1.64u w=0.265u l=0.28u
X1 S_uq0 a_136_n44# D VSUBS nfet_03v3 ad=0.15742p pd=1.65u as=91.3f ps=0.92u w=0.265u l=0.28u
.ends

.subckt ypass_gate_a_3v1024x8m81 b bb ypass pcb vdd_uq0 m3_n41_6881# m3_n41_5924#
+ m3_n41_6639# vss m3_n41_4610# m3_n41_5682# m3_n41_6398# vdd pmos_5p0431059130201_3v1024x8m81_0/D
+ pmos_5p0431059130201_3v1024x8m81_1/D pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ m3_n41_5198# m3_n41_5440# m3_n41_6156#
Xpmos_1p2$$46889004_3v1024x8m81_1 pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ nmos_5p0431059130202_3v1024x8m81_0/D vdd_uq0 pmos_5p0431059130201_3v1024x8m81_0/D
+ pmos_1p2$$46889004_3v1024x8m81
Xnmos_1p2$$47119404_3v1024x8m81_1 pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass pmos_5p0431059130201_3v1024x8m81_0/D vss nmos_1p2$$47119404_3v1024x8m81
Xpmos_5p0431059130201_3v1024x8m81_0 pmos_5p0431059130201_3v1024x8m81_0/D pcb vdd bb
+ pmos_5p0431059130201_3v1024x8m81
Xnmos_1p2$$47119404_3v1024x8m81_3 pmos_5p0431059130201_3v1024x8m81_1/D ypass bb vss
+ nmos_1p2$$47119404_3v1024x8m81
Xpmos_5p0431059130201_3v1024x8m81_1 pmos_5p0431059130201_3v1024x8m81_1/D nmos_5p0431059130202_3v1024x8m81_0/D
+ vdd bb pmos_5p0431059130201_3v1024x8m81
Xnmos_5p0431059130202_3v1024x8m81_0 nmos_5p0431059130202_3v1024x8m81_0/D ypass ypass
+ vss vss vss nmos_5p0431059130202_3v1024x8m81
X0 vdd pcb pmos_5p0431059130201_3v1024x8m81_0/D vdd pfet_03v3 ad=1.06988p pd=4.52u as=0.4121p ps=2.105u w=1.585u l=0.28u
X1 pmos_5p0431059130201_3v1024x8m81_0/D pcb vdd vdd pfet_03v3 ad=0.4121p pd=2.105u as=0.99855p ps=4.43u w=1.585u l=0.28u
X2 vdd_uq0 ypass nmos_5p0431059130202_3v1024x8m81_0/D vdd_uq0 pfet_03v3 ad=0.5143p pd=2.87u as=0.34055p ps=1.675u w=0.695u l=0.28u
X3 vdd pcb bb vdd pfet_03v3 ad=1.07325p pd=4.53u as=0.4134p ps=2.11u w=1.59u l=0.28u
X4 bb pcb vdd vdd pfet_03v3 ad=0.4134p pd=2.11u as=1.0017p ps=4.44u w=1.59u l=0.28u
X5 nmos_5p0431059130202_3v1024x8m81_0/D ypass vdd_uq0 vdd_uq0 pfet_03v3 ad=0.34055p pd=1.675u as=0.38572p ps=2.5u w=0.695u l=0.28u
.ends

.subckt ypass_gate_3v1024x8m81 vdd b bb ypass pcb vdd_uq0 m3_n41_6881# m3_n41_5924#
+ m3_n41_6639# m3_n41_4610# pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ m3_n41_5682# m3_n41_6398# db m3_n41_5198# m3_n41_5440# m3_n41_6156# vss
Xpmos_1p2$$46889004_3v1024x8m81_1 pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ nmos_5p0431059130202_3v1024x8m81_0/D vdd_uq0 b pmos_1p2$$46889004_3v1024x8m81
Xnmos_1p2$$47119404_3v1024x8m81_1 pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass b vss nmos_1p2$$47119404_3v1024x8m81
Xpmos_5p0431059130201_3v1024x8m81_0 b pcb vdd bb pmos_5p0431059130201_3v1024x8m81
Xnmos_1p2$$47119404_3v1024x8m81_3 db ypass bb vss nmos_1p2$$47119404_3v1024x8m81
Xpmos_5p0431059130201_3v1024x8m81_1 db nmos_5p0431059130202_3v1024x8m81_0/D vdd bb
+ pmos_5p0431059130201_3v1024x8m81
Xnmos_5p0431059130202_3v1024x8m81_0 nmos_5p0431059130202_3v1024x8m81_0/D ypass ypass
+ vss vss vss nmos_5p0431059130202_3v1024x8m81
X0 vdd pcb b vdd pfet_03v3 ad=0.92722p pd=4.34u as=0.4121p ps=2.105u w=1.585u l=0.28u
X1 b pcb vdd vdd pfet_03v3 ad=0.4121p pd=2.105u as=0.93515p ps=4.35u w=1.585u l=0.28u
X2 nmos_5p0431059130202_3v1024x8m81_0/D ypass vdd_uq0 vdd_uq0 pfet_03v3 ad=0.26235p pd=1.45u as=0.46218p ps=2.72u w=0.695u l=0.28u
X3 vdd_uq0 ypass nmos_5p0431059130202_3v1024x8m81_0/D vdd_uq0 pfet_03v3 ad=0.39963p pd=2.54u as=0.26235p ps=1.45u w=0.695u l=0.28u
X4 vdd pcb bb vdd pfet_03v3 ad=0.93015p pd=4.35u as=0.4134p ps=2.11u w=1.59u l=0.28u
X5 bb pcb vdd vdd pfet_03v3 ad=0.4134p pd=2.11u as=0.9381p ps=4.36u w=1.59u l=0.28u
.ends

.subckt mux821_3v1024x8m81 ypass_gate_3v1024x8m81_6/b ypass_gate_3v1024x8m81_6/bb
+ ypass_gate_3v1024x8m81_3/bb ypass_gate_3v1024x8m81_7/db ypass_gate_3v1024x8m81_6/pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_5/db ypass_gate_a_3v1024x8m81_0/ypass ypass_gate_3v1024x8m81_1/b
+ ypass_gate_3v1024x8m81_1/ypass ypass_gate_3v1024x8m81_2/ypass ypass_gate_a_3v1024x8m81_0/bb
+ ypass_gate_3v1024x8m81_5/bb ypass_gate_3v1024x8m81_3/ypass ypass_gate_3v1024x8m81_4/pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_3/b ypass_gate_3v1024x8m81_2/bb ypass_gate_3v1024x8m81_4/ypass
+ ypass_gate_3v1024x8m81_5/ypass ypass_gate_3v1024x8m81_5/b ypass_gate_3v1024x8m81_6/ypass
+ ypass_gate_3v1024x8m81_7/pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_7/ypass ypass_gate_3v1024x8m81_7/b ypass_gate_a_3v1024x8m81_0/pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_7/bb ypass_gate_3v1024x8m81_5/pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_4/bb ypass_gate_3v1024x8m81_1/bb ypass_gate_3v1024x8m81_4/db
+ ypass_gate_3v1024x8m81_1/db ypass_gate_3v1024x8m81_2/pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_7/m3_n41_5924# ypass_gate_3v1024x8m81_7/m3_n41_6881# ypass_gate_3v1024x8m81_7/m3_n41_5682#
+ ypass_gate_3v1024x8m81_7/m3_n41_5198# ypass_gate_3v1024x8m81_2/b ypass_gate_3v1024x8m81_7/vdd_uq0
+ ypass_gate_3v1024x8m81_7/m3_n41_6398# ypass_gate_3v1024x8m81_7/m3_n41_5440# ypass_gate_3v1024x8m81_7/m3_n41_6156#
+ ypass_gate_3v1024x8m81_3/pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_a_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D ypass_gate_3v1024x8m81_4/b
+ ypass_gate_3v1024x8m81_7/vdd VSUBS ypass_gate_3v1024x8m81_7/m3_n41_6639# ypass_gate_3v1024x8m81_1/pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_7/pcb
Xypass_gate_a_3v1024x8m81_0 ypass_gate_a_3v1024x8m81_0/b ypass_gate_a_3v1024x8m81_0/bb
+ ypass_gate_a_3v1024x8m81_0/ypass ypass_gate_3v1024x8m81_7/pcb ypass_gate_3v1024x8m81_7/vdd_uq0
+ ypass_gate_3v1024x8m81_7/m3_n41_6881# ypass_gate_3v1024x8m81_7/m3_n41_5924# ypass_gate_3v1024x8m81_7/m3_n41_6639#
+ VSUBS ypass_gate_3v1024x8m81_7/vdd_uq0 ypass_gate_3v1024x8m81_7/m3_n41_5682# ypass_gate_3v1024x8m81_7/m3_n41_6398#
+ ypass_gate_3v1024x8m81_7/vdd ypass_gate_a_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_1/db ypass_gate_a_3v1024x8m81_0/pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_7/m3_n41_5198# ypass_gate_3v1024x8m81_7/m3_n41_5440# ypass_gate_3v1024x8m81_7/m3_n41_6156#
+ ypass_gate_a_3v1024x8m81
Xypass_gate_3v1024x8m81_1 ypass_gate_3v1024x8m81_7/vdd ypass_gate_3v1024x8m81_1/b
+ ypass_gate_3v1024x8m81_1/bb ypass_gate_3v1024x8m81_1/ypass ypass_gate_3v1024x8m81_7/pcb
+ ypass_gate_3v1024x8m81_7/vdd_uq0 ypass_gate_3v1024x8m81_7/m3_n41_6881# ypass_gate_3v1024x8m81_7/m3_n41_5924#
+ ypass_gate_3v1024x8m81_7/m3_n41_6639# ypass_gate_3v1024x8m81_7/vdd_uq0 ypass_gate_3v1024x8m81_1/pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_7/m3_n41_5682# ypass_gate_3v1024x8m81_7/m3_n41_6398# ypass_gate_3v1024x8m81_1/db
+ ypass_gate_3v1024x8m81_7/m3_n41_5198# ypass_gate_3v1024x8m81_7/m3_n41_5440# ypass_gate_3v1024x8m81_7/m3_n41_6156#
+ VSUBS ypass_gate_3v1024x8m81
Xypass_gate_3v1024x8m81_2 ypass_gate_3v1024x8m81_7/vdd ypass_gate_3v1024x8m81_2/b
+ ypass_gate_3v1024x8m81_2/bb ypass_gate_3v1024x8m81_2/ypass ypass_gate_3v1024x8m81_7/pcb
+ ypass_gate_3v1024x8m81_7/vdd_uq0 ypass_gate_3v1024x8m81_7/m3_n41_6881# ypass_gate_3v1024x8m81_7/m3_n41_5924#
+ ypass_gate_3v1024x8m81_7/m3_n41_6639# ypass_gate_3v1024x8m81_7/vdd_uq0 ypass_gate_3v1024x8m81_2/pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_7/m3_n41_5682# ypass_gate_3v1024x8m81_7/m3_n41_6398# ypass_gate_3v1024x8m81_4/db
+ ypass_gate_3v1024x8m81_7/m3_n41_5198# ypass_gate_3v1024x8m81_7/m3_n41_5440# ypass_gate_3v1024x8m81_7/m3_n41_6156#
+ VSUBS ypass_gate_3v1024x8m81
Xypass_gate_3v1024x8m81_3 ypass_gate_3v1024x8m81_7/vdd ypass_gate_3v1024x8m81_3/b
+ ypass_gate_3v1024x8m81_3/bb ypass_gate_3v1024x8m81_3/ypass ypass_gate_3v1024x8m81_7/pcb
+ ypass_gate_3v1024x8m81_7/vdd_uq0 ypass_gate_3v1024x8m81_7/m3_n41_6881# ypass_gate_3v1024x8m81_7/m3_n41_5924#
+ ypass_gate_3v1024x8m81_7/m3_n41_6639# ypass_gate_3v1024x8m81_7/vdd_uq0 ypass_gate_3v1024x8m81_3/pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_7/m3_n41_5682# ypass_gate_3v1024x8m81_7/m3_n41_6398# ypass_gate_3v1024x8m81_5/db
+ ypass_gate_3v1024x8m81_7/m3_n41_5198# ypass_gate_3v1024x8m81_7/m3_n41_5440# ypass_gate_3v1024x8m81_7/m3_n41_6156#
+ VSUBS ypass_gate_3v1024x8m81
Xypass_gate_3v1024x8m81_4 ypass_gate_3v1024x8m81_7/vdd ypass_gate_3v1024x8m81_4/b
+ ypass_gate_3v1024x8m81_4/bb ypass_gate_3v1024x8m81_4/ypass ypass_gate_3v1024x8m81_7/pcb
+ ypass_gate_3v1024x8m81_7/vdd_uq0 ypass_gate_3v1024x8m81_7/m3_n41_6881# ypass_gate_3v1024x8m81_7/m3_n41_5924#
+ ypass_gate_3v1024x8m81_7/m3_n41_6639# ypass_gate_3v1024x8m81_7/vdd_uq0 ypass_gate_3v1024x8m81_4/pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_7/m3_n41_5682# ypass_gate_3v1024x8m81_7/m3_n41_6398# ypass_gate_3v1024x8m81_4/db
+ ypass_gate_3v1024x8m81_7/m3_n41_5198# ypass_gate_3v1024x8m81_7/m3_n41_5440# ypass_gate_3v1024x8m81_7/m3_n41_6156#
+ VSUBS ypass_gate_3v1024x8m81
Xypass_gate_3v1024x8m81_5 ypass_gate_3v1024x8m81_7/vdd ypass_gate_3v1024x8m81_5/b
+ ypass_gate_3v1024x8m81_5/bb ypass_gate_3v1024x8m81_5/ypass ypass_gate_3v1024x8m81_7/pcb
+ ypass_gate_3v1024x8m81_7/vdd_uq0 ypass_gate_3v1024x8m81_7/m3_n41_6881# ypass_gate_3v1024x8m81_7/m3_n41_5924#
+ ypass_gate_3v1024x8m81_7/m3_n41_6639# ypass_gate_3v1024x8m81_7/vdd_uq0 ypass_gate_3v1024x8m81_5/pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_7/m3_n41_5682# ypass_gate_3v1024x8m81_7/m3_n41_6398# ypass_gate_3v1024x8m81_5/db
+ ypass_gate_3v1024x8m81_7/m3_n41_5198# ypass_gate_3v1024x8m81_7/m3_n41_5440# ypass_gate_3v1024x8m81_7/m3_n41_6156#
+ VSUBS ypass_gate_3v1024x8m81
Xypass_gate_3v1024x8m81_6 ypass_gate_3v1024x8m81_7/vdd ypass_gate_3v1024x8m81_6/b
+ ypass_gate_3v1024x8m81_6/bb ypass_gate_3v1024x8m81_6/ypass ypass_gate_3v1024x8m81_7/pcb
+ ypass_gate_3v1024x8m81_7/vdd_uq0 ypass_gate_3v1024x8m81_7/m3_n41_6881# ypass_gate_3v1024x8m81_7/m3_n41_5924#
+ ypass_gate_3v1024x8m81_7/m3_n41_6639# ypass_gate_3v1024x8m81_7/vdd_uq0 ypass_gate_3v1024x8m81_6/pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_7/m3_n41_5682# ypass_gate_3v1024x8m81_7/m3_n41_6398# ypass_gate_3v1024x8m81_7/db
+ ypass_gate_3v1024x8m81_7/m3_n41_5198# ypass_gate_3v1024x8m81_7/m3_n41_5440# ypass_gate_3v1024x8m81_7/m3_n41_6156#
+ VSUBS ypass_gate_3v1024x8m81
Xypass_gate_3v1024x8m81_7 ypass_gate_3v1024x8m81_7/vdd ypass_gate_3v1024x8m81_7/b
+ ypass_gate_3v1024x8m81_7/bb ypass_gate_3v1024x8m81_7/ypass ypass_gate_3v1024x8m81_7/pcb
+ ypass_gate_3v1024x8m81_7/vdd_uq0 ypass_gate_3v1024x8m81_7/m3_n41_6881# ypass_gate_3v1024x8m81_7/m3_n41_5924#
+ ypass_gate_3v1024x8m81_7/m3_n41_6639# ypass_gate_3v1024x8m81_7/vdd_uq0 ypass_gate_3v1024x8m81_7/pmos_1p2$$46889004_3v1024x8m81_1/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_7/m3_n41_5682# ypass_gate_3v1024x8m81_7/m3_n41_6398# ypass_gate_3v1024x8m81_7/db
+ ypass_gate_3v1024x8m81_7/m3_n41_5198# ypass_gate_3v1024x8m81_7/m3_n41_5440# ypass_gate_3v1024x8m81_7/m3_n41_6156#
+ VSUBS ypass_gate_3v1024x8m81
.ends

.subckt pmos_1p2$$202583084_3v1024x8m81 a_n42_n34# w_n133_n66# pmos_5p04310591302035_3v1024x8m81_0/S_uq0
+ pmos_5p04310591302035_3v1024x8m81_0/S a_118_n34# pmos_5p04310591302035_3v1024x8m81_0/D
Xpmos_5p04310591302035_3v1024x8m81_0 pmos_5p04310591302035_3v1024x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302035_3v1024x8m81_0/S_uq0 pmos_5p04310591302035_3v1024x8m81_0/S
+ pmos_5p04310591302035_3v1024x8m81
.ends

.subckt nmos_5p04310591302040_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.2794p pd=2.15u as=0.2794p ps=2.15u w=0.635u l=0.28u
.ends

.subckt pmos_1p2$$202585132_3v1024x8m81 a_n14_n34# pmos_5p04310591302014_3v1024x8m81_0/S
+ w_n119_n65# pmos_5p04310591302014_3v1024x8m81_0/D
Xpmos_5p04310591302014_3v1024x8m81_0 pmos_5p04310591302014_3v1024x8m81_0/D a_n14_n34#
+ w_n119_n65# pmos_5p04310591302014_3v1024x8m81_0/S pmos_5p04310591302014_3v1024x8m81
.ends

.subckt pmos_5p04310591302043_3v1024x8m81 D_uq0 D a_265_n44# S_uq0 S a_n56_n44# a_104_n44#
+ w_n230_n86#
X0 D_uq0 a_265_n44# S_uq0 w_n230_n86# pfet_03v3 ad=0.4092p pd=2.74u as=0.24412p ps=1.455u w=0.93u l=0.28u
X1 D a_n56_n44# S w_n230_n86# pfet_03v3 ad=0.2418p pd=1.45u as=0.4092p ps=2.74u w=0.93u l=0.28u
X2 S_uq0 a_104_n44# D w_n230_n86# pfet_03v3 ad=0.24412p pd=1.455u as=0.2418p ps=1.45u w=0.93u l=0.28u
.ends

.subckt nmos_1p2$$202595372_3v1024x8m81 nmos_5p0431059130208_3v1024x8m81_0/S nmos_5p0431059130208_3v1024x8m81_0/D
+ a_n14_89# VSUBS
Xnmos_5p0431059130208_3v1024x8m81_0 nmos_5p0431059130208_3v1024x8m81_0/D a_n14_89#
+ nmos_5p0431059130208_3v1024x8m81_0/S VSUBS nmos_5p0431059130208_3v1024x8m81
.ends

.subckt pmos_1p2$$202584108_3v1024x8m81 a_n14_n34# pmos_5p04310591302014_3v1024x8m81_0/S
+ pmos_5p04310591302014_3v1024x8m81_0/D w_n133_n65#
Xpmos_5p04310591302014_3v1024x8m81_0 pmos_5p04310591302014_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302014_3v1024x8m81_0/S pmos_5p04310591302014_3v1024x8m81
.ends

.subckt pmos_1p2$$202587180_3v1024x8m81 a_n14_n34# pmos_5p04310591302014_3v1024x8m81_0/S
+ pmos_5p04310591302014_3v1024x8m81_0/D w_n133_n65#
Xpmos_5p04310591302014_3v1024x8m81_0 pmos_5p04310591302014_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302014_3v1024x8m81_0/S pmos_5p04310591302014_3v1024x8m81
.ends

.subckt nmos_5p04310591302042_3v1024x8m81 D_uq0 D a_265_n44# S_uq0 S a_n56_n44# a_104_n44#
+ VSUBS
X0 D_uq0 a_265_n44# S_uq0 VSUBS nfet_03v3 ad=0.1628p pd=1.62u as=97.125f ps=0.895u w=0.37u l=0.28u
X1 D a_n56_n44# S VSUBS nfet_03v3 ad=96.2f pd=0.89u as=0.1628p ps=1.62u w=0.37u l=0.28u
X2 S_uq0 a_104_n44# D VSUBS nfet_03v3 ad=97.125f pd=0.895u as=96.2f ps=0.89u w=0.37u l=0.28u
.ends

.subckt nmos_1p2$$202594348_3v1024x8m81 nmos_5p04310591302040_3v1024x8m81_0/D nmos_5p04310591302040_3v1024x8m81_0/S
+ a_n14_n44# VSUBS
Xnmos_5p04310591302040_3v1024x8m81_0 nmos_5p04310591302040_3v1024x8m81_0/D a_n14_n44#
+ nmos_5p04310591302040_3v1024x8m81_0/S VSUBS nmos_5p04310591302040_3v1024x8m81
.ends

.subckt pmos_1p2$$202586156_3v1024x8m81 a_n14_n34# pmos_5p04310591302014_3v1024x8m81_0/S
+ pmos_5p04310591302014_3v1024x8m81_0/D w_n133_n65#
Xpmos_5p04310591302014_3v1024x8m81_0 pmos_5p04310591302014_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302014_3v1024x8m81_0/S pmos_5p04310591302014_3v1024x8m81
.ends

.subckt nmos_1p2$$202596396_3v1024x8m81 nmos_5p0431059130208_3v1024x8m81_0/S nmos_5p0431059130208_3v1024x8m81_0/D
+ a_n14_89# VSUBS
Xnmos_5p0431059130208_3v1024x8m81_0 nmos_5p0431059130208_3v1024x8m81_0/D a_n14_89#
+ nmos_5p0431059130208_3v1024x8m81_0/S VSUBS nmos_5p0431059130208_3v1024x8m81
.ends

.subckt nmos_1p2$$202598444_3v1024x8m81 nmos_5p04310591302010_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v1024x8m81_0/S VSUBS
Xnmos_5p04310591302010_3v1024x8m81_0 nmos_5p04310591302010_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v1024x8m81_0/S VSUBS nmos_5p04310591302010_3v1024x8m81
.ends

.subckt pmos_5p04310591302041_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
.ends

.subckt nmos_5p04310591302039_3v1024x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt wen_wm1_3v1024x8m81 GWEN men wep vdd wen vss vdd_uq0
Xpmos_1p2$$202583084_3v1024x8m81_0 nmos_1p2$$202596396_3v1024x8m81_0/nmos_5p0431059130208_3v1024x8m81_0/D
+ vdd vdd vdd nmos_1p2$$202596396_3v1024x8m81_0/nmos_5p0431059130208_3v1024x8m81_0/D
+ pmos_1p2$$202583084_3v1024x8m81_0/pmos_5p04310591302035_3v1024x8m81_0/D pmos_1p2$$202583084_3v1024x8m81
Xnmos_5p04310591302040_3v1024x8m81_0 pmos_5p04310591302035_3v1024x8m81_0/D pmos_5p04310591302020_3v1024x8m81_0/S
+ vss vss nmos_5p04310591302040_3v1024x8m81
Xnmos_5p04310591302040_3v1024x8m81_1 pmos_5p04310591302014_3v1024x8m81_5/D men vss
+ vss nmos_5p04310591302040_3v1024x8m81
Xpmos_1p2$$202585132_3v1024x8m81_0 nmos_1p2$$202595372_3v1024x8m81_1/nmos_5p0431059130208_3v1024x8m81_0/S
+ vdd vdd nmos_1p2$$202596396_3v1024x8m81_0/nmos_5p0431059130208_3v1024x8m81_0/D pmos_1p2$$202585132_3v1024x8m81
Xnmos_5p04310591302040_3v1024x8m81_2 vss vss pmos_5p04310591302014_3v1024x8m81_5/D
+ vss nmos_5p04310591302040_3v1024x8m81
Xpmos_5p04310591302043_3v1024x8m81_0 wep wep pmos_5p04310591302035_3v1024x8m81_0/D
+ vdd_uq0 vdd_uq0 pmos_5p04310591302035_3v1024x8m81_0/D pmos_5p04310591302035_3v1024x8m81_0/D
+ vdd_uq0 pmos_5p04310591302043_3v1024x8m81
Xnmos_5p0431059130208_3v1024x8m81_0 vss GWEN nmos_5p0431059130208_3v1024x8m81_2/D
+ vss nmos_5p0431059130208_3v1024x8m81
Xnmos_5p0431059130208_3v1024x8m81_1 nmos_5p0431059130208_3v1024x8m81_1/D nmos_5p0431059130208_3v1024x8m81_2/D
+ vss vss nmos_5p0431059130208_3v1024x8m81
Xnmos_1p2$$202595372_3v1024x8m81_0 pmos_5p04310591302041_3v1024x8m81_0/S pmos_5p04310591302041_3v1024x8m81_0/D
+ nmos_5p0431059130208_3v1024x8m81_3/D vss nmos_1p2$$202595372_3v1024x8m81
Xpmos_1p2$$202584108_3v1024x8m81_0 pmos_5p04310591302041_3v1024x8m81_0/S nmos_1p2$$202595372_3v1024x8m81_1/nmos_5p0431059130208_3v1024x8m81_0/S
+ vdd vdd pmos_1p2$$202584108_3v1024x8m81
Xnmos_5p0431059130208_3v1024x8m81_2 nmos_5p0431059130208_3v1024x8m81_2/D wen vss vss
+ nmos_5p0431059130208_3v1024x8m81
Xnmos_1p2$$202595372_3v1024x8m81_1 nmos_1p2$$202595372_3v1024x8m81_1/nmos_5p0431059130208_3v1024x8m81_0/S
+ vss pmos_5p04310591302041_3v1024x8m81_0/S vss nmos_1p2$$202595372_3v1024x8m81
Xnmos_5p0431059130208_3v1024x8m81_3 nmos_5p0431059130208_3v1024x8m81_3/D pmos_5p04310591302014_3v1024x8m81_5/D
+ vss vss nmos_5p0431059130208_3v1024x8m81
Xpmos_1p2$$202587180_3v1024x8m81_0 nmos_5p0431059130208_3v1024x8m81_3/D nmos_5p0431059130208_3v1024x8m81_1/D
+ pmos_5p04310591302041_3v1024x8m81_0/S vdd pmos_1p2$$202587180_3v1024x8m81
Xnmos_5p04310591302042_3v1024x8m81_0 wep wep pmos_5p04310591302035_3v1024x8m81_0/D
+ vss vss pmos_5p04310591302035_3v1024x8m81_0/D pmos_5p04310591302035_3v1024x8m81_0/D
+ vss nmos_5p04310591302042_3v1024x8m81
Xnmos_1p2$$202594348_3v1024x8m81_0 vss pmos_1p2$$202583084_3v1024x8m81_0/pmos_5p04310591302035_3v1024x8m81_0/D
+ nmos_1p2$$202596396_3v1024x8m81_0/nmos_5p0431059130208_3v1024x8m81_0/D vss nmos_1p2$$202594348_3v1024x8m81
Xpmos_1p2$$202586156_3v1024x8m81_0 nmos_1p2$$202595372_3v1024x8m81_1/nmos_5p0431059130208_3v1024x8m81_0/S
+ pmos_5p04310591302041_3v1024x8m81_0/D vdd vdd pmos_1p2$$202586156_3v1024x8m81
Xpmos_5p04310591302014_3v1024x8m81_0 pmos_5p04310591302014_3v1024x8m81_2/S wen vdd_uq0
+ vdd_uq0 pmos_5p04310591302014_3v1024x8m81
Xpmos_5p04310591302014_3v1024x8m81_1 nmos_5p0431059130208_3v1024x8m81_1/D nmos_5p0431059130208_3v1024x8m81_2/D
+ vdd_uq0 vdd_uq0 pmos_5p04310591302014_3v1024x8m81
Xpmos_5p04310591302014_3v1024x8m81_2 nmos_5p0431059130208_3v1024x8m81_2/D GWEN vdd_uq0
+ pmos_5p04310591302014_3v1024x8m81_2/S pmos_5p04310591302014_3v1024x8m81
Xnmos_1p2$$202596396_3v1024x8m81_0 vss nmos_1p2$$202596396_3v1024x8m81_0/nmos_5p0431059130208_3v1024x8m81_0/D
+ nmos_1p2$$202595372_3v1024x8m81_1/nmos_5p0431059130208_3v1024x8m81_0/S vss nmos_1p2$$202596396_3v1024x8m81
Xpmos_5p04310591302014_3v1024x8m81_3 pmos_5p04310591302014_3v1024x8m81_5/S men vdd
+ vdd pmos_5p04310591302014_3v1024x8m81
Xpmos_5p04310591302035_3v1024x8m81_0 pmos_5p04310591302035_3v1024x8m81_0/D pmos_5p04310591302020_3v1024x8m81_0/S
+ pmos_5p04310591302020_3v1024x8m81_0/S vdd_uq0 vdd_uq0 vdd_uq0 pmos_5p04310591302035_3v1024x8m81
Xnmos_1p2$$202596396_3v1024x8m81_1 pmos_5p04310591302041_3v1024x8m81_0/D vss nmos_1p2$$202595372_3v1024x8m81_1/nmos_5p0431059130208_3v1024x8m81_0/S
+ vss nmos_1p2$$202596396_3v1024x8m81
Xpmos_5p04310591302014_3v1024x8m81_4 nmos_5p0431059130208_3v1024x8m81_3/D pmos_5p04310591302014_3v1024x8m81_5/D
+ vdd vdd pmos_5p04310591302014_3v1024x8m81
Xpmos_5p04310591302014_3v1024x8m81_5 pmos_5p04310591302014_3v1024x8m81_5/D vss vdd
+ pmos_5p04310591302014_3v1024x8m81_5/S pmos_5p04310591302014_3v1024x8m81
Xnmos_1p2$$202598444_3v1024x8m81_0 pmos_5p04310591302041_3v1024x8m81_0/S pmos_5p04310591302014_3v1024x8m81_5/D
+ nmos_5p0431059130208_3v1024x8m81_1/D vss nmos_1p2$$202598444_3v1024x8m81
Xpmos_5p04310591302020_3v1024x8m81_0 men nmos_1p2$$202596396_3v1024x8m81_0/nmos_5p0431059130208_3v1024x8m81_0/D
+ nmos_1p2$$202596396_3v1024x8m81_0/nmos_5p0431059130208_3v1024x8m81_0/D vdd pmos_5p04310591302020_3v1024x8m81_0/S
+ pmos_5p04310591302020_3v1024x8m81_0/S pmos_5p04310591302020_3v1024x8m81
Xnmos_5p04310591302010_3v1024x8m81_0 vss nmos_1p2$$202596396_3v1024x8m81_0/nmos_5p0431059130208_3v1024x8m81_0/D
+ pmos_5p04310591302020_3v1024x8m81_0/S vss nmos_5p04310591302010_3v1024x8m81
Xpmos_5p04310591302041_3v1024x8m81_0 pmos_5p04310591302041_3v1024x8m81_0/D pmos_5p04310591302014_3v1024x8m81_5/D
+ vdd pmos_5p04310591302041_3v1024x8m81_0/S pmos_5p04310591302041_3v1024x8m81
Xnmos_5p04310591302039_3v1024x8m81_0 men pmos_1p2$$202583084_3v1024x8m81_0/pmos_5p04310591302035_3v1024x8m81_0/D
+ pmos_1p2$$202583084_3v1024x8m81_0/pmos_5p04310591302035_3v1024x8m81_0/D pmos_5p04310591302020_3v1024x8m81_0/S
+ pmos_5p04310591302020_3v1024x8m81_0/S vss nmos_5p04310591302039_3v1024x8m81
.ends

.subckt nmos_5p04310591302052_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.3278p pd=2.37u as=0.3278p ps=2.37u w=0.745u l=0.28u
.ends

.subckt nmos_5p04310591302045_3v1024x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.583p ps=3.53u w=1.325u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.583p pd=3.53u as=0.3445p ps=1.845u w=1.325u l=0.28u
.ends

.subckt pmos_5p04310591302048_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.924p pd=5.08u as=0.924p ps=5.08u w=2.1u l=0.28u
.ends

.subckt nmos_5p04310591302044_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.451p pd=2.93u as=0.451p ps=2.93u w=1.025u l=0.28u
.ends

.subckt pmos_5p04310591302051_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.6877p pd=3.165u as=1.1638p ps=6.17u w=2.645u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=1.1638p pd=6.17u as=0.6877p ps=3.165u w=2.645u l=0.28u
.ends

.subckt pmos_5p04310591302047_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.8206p pd=4.61u as=0.8206p ps=4.61u w=1.865u l=0.28u
.ends

.subckt nmos_5p04310591302050_3v1024x8m81 D_uq0 D a_265_n44# S_uq0 S a_n56_n44# a_104_n44#
+ VSUBS
X0 D_uq0 a_265_n44# S_uq0 VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.27692p ps=1.58u w=1.055u l=0.28u
X1 D a_n56_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X2 S_uq0 a_104_n44# D VSUBS nfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt nmos_5p04310591302046_3v1024x8m81 a_20_n44# D_uq1 D_uq0 D a_181_n44# a_502_n44#
+ S_uq2 a_662_n44# S_uq1 a_n140_n44# S_uq0 S a_341_n44# VSUBS
X0 S a_341_n44# D VSUBS nfet_03v3 ad=0.25855p pd=1.51u as=0.2561p ps=1.505u w=0.985u l=0.28u
X1 S_uq0 a_662_n44# D_uq0 VSUBS nfet_03v3 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.28u
X2 D_uq0 a_502_n44# S VSUBS nfet_03v3 ad=0.2561p pd=1.505u as=0.25855p ps=1.51u w=0.985u l=0.28u
X3 S_uq1 a_20_n44# D_uq1 VSUBS nfet_03v3 ad=0.25855p pd=1.51u as=0.2561p ps=1.505u w=0.985u l=0.28u
X4 D a_181_n44# S_uq1 VSUBS nfet_03v3 ad=0.2561p pd=1.505u as=0.25855p ps=1.51u w=0.985u l=0.28u
X5 D_uq1 a_n140_n44# S_uq2 VSUBS nfet_03v3 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.28u
.ends

.subckt pmos_5p04310591302049_3v1024x8m81 a_20_n44# D_uq1 D_uq0 D a_181_n44# S_uq2
+ S_uq1 a_n140_n44# S_uq0 S a_341_n44# a_503_n44# a_663_n44# w_n314_n86#
X0 S a_341_n44# D w_n314_n86# pfet_03v3 ad=0.4664p pd=2.29u as=0.4576p ps=2.28u w=1.76u l=0.28u
X1 S_uq1 a_20_n44# D_uq1 w_n314_n86# pfet_03v3 ad=0.462p pd=2.285u as=0.4576p ps=2.28u w=1.76u l=0.28u
X2 D a_181_n44# S_uq1 w_n314_n86# pfet_03v3 ad=0.4576p pd=2.28u as=0.462p ps=2.285u w=1.76u l=0.28u
X3 D_uq1 a_n140_n44# S_uq2 w_n314_n86# pfet_03v3 ad=0.4576p pd=2.28u as=0.7744p ps=4.4u w=1.76u l=0.28u
X4 S_uq0 a_663_n44# D_uq0 w_n314_n86# pfet_03v3 ad=0.7832p pd=4.41u as=0.4576p ps=2.28u w=1.76u l=0.28u
X5 D_uq0 a_503_n44# S w_n314_n86# pfet_03v3 ad=0.4576p pd=2.28u as=0.4664p ps=2.29u w=1.76u l=0.28u
.ends

.subckt pmos_1p2$$171625516_3v1024x8m81 a_n42_n34# pmos_5p0431059130203_3v1024x8m81_0/w_n202_n86#
+ pmos_5p0431059130203_3v1024x8m81_0/S a_118_n34# pmos_5p0431059130203_3v1024x8m81_0/D
+ pmos_5p0431059130203_3v1024x8m81_0/S_uq0
Xpmos_5p0431059130203_3v1024x8m81_0 pmos_5p0431059130203_3v1024x8m81_0/D a_n42_n34#
+ a_118_n34# pmos_5p0431059130203_3v1024x8m81_0/w_n202_n86# pmos_5p0431059130203_3v1024x8m81_0/S_uq0
+ pmos_5p0431059130203_3v1024x8m81_0/S pmos_5p0431059130203_3v1024x8m81
.ends

.subckt outbuf_oe_3v1024x8m81 qp qn se q GWE vss vdd
Xnmos_5p04310591302052_3v1024x8m81_0 vss GWE pmos_5p04310591302047_3v1024x8m81_0/S
+ vss nmos_5p04310591302052_3v1024x8m81
Xnmos_5p04310591302045_3v1024x8m81_0 vss pmos_5p04310591302047_3v1024x8m81_0/S pmos_5p04310591302047_3v1024x8m81_0/S
+ nmos_5p04310591302045_3v1024x8m81_1/S nmos_5p04310591302045_3v1024x8m81_1/S vss
+ nmos_5p04310591302045_3v1024x8m81
Xnmos_5p0431059130208_3v1024x8m81_0 nmos_5p0431059130208_3v1024x8m81_0/D se vss vss
+ nmos_5p0431059130208_3v1024x8m81
Xnmos_5p04310591302033_3v1024x8m81_0 pmos_5p04310591302038_3v1024x8m81_0/D pmos_5p04310591302051_3v1024x8m81_0/D
+ vss vss nmos_5p04310591302033_3v1024x8m81
Xnmos_5p04310591302045_3v1024x8m81_1 pmos_5p04310591302051_3v1024x8m81_0/D qn qn nmos_5p04310591302045_3v1024x8m81_1/S
+ nmos_5p04310591302045_3v1024x8m81_1/S vss nmos_5p04310591302045_3v1024x8m81
Xnmos_5p0431059130208_3v1024x8m81_1 vss pmos_5p04310591302038_3v1024x8m81_0/D nmos_5p0431059130208_3v1024x8m81_1/S
+ vss nmos_5p0431059130208_3v1024x8m81
Xpmos_5p04310591302048_3v1024x8m81_0 vdd pmos_5p04310591302047_3v1024x8m81_0/S vdd
+ pmos_5p04310591302048_3v1024x8m81_0/S pmos_5p04310591302048_3v1024x8m81
Xnmos_5p04310591302044_3v1024x8m81_0 vss pmos_5p04310591302047_3v1024x8m81_0/S pmos_5p04310591302048_3v1024x8m81_0/S
+ vss nmos_5p04310591302044_3v1024x8m81
Xpmos_5p04310591302014_3v1024x8m81_0 nmos_5p0431059130208_3v1024x8m81_0/D se vdd vdd
+ pmos_5p04310591302014_3v1024x8m81
Xpmos_5p04310591302038_3v1024x8m81_0 pmos_5p04310591302038_3v1024x8m81_0/D pmos_5p04310591302051_3v1024x8m81_0/D
+ vdd vdd pmos_5p04310591302038_3v1024x8m81
Xpmos_5p04310591302051_3v1024x8m81_0 pmos_5p04310591302051_3v1024x8m81_0/D qp qp vdd
+ pmos_5p04310591302051_3v1024x8m81_1/S pmos_5p04310591302051_3v1024x8m81_1/S pmos_5p04310591302051_3v1024x8m81
Xpmos_5p04310591302047_3v1024x8m81_0 vdd GWE vdd pmos_5p04310591302047_3v1024x8m81_0/S
+ pmos_5p04310591302047_3v1024x8m81
Xpmos_5p04310591302051_3v1024x8m81_1 vdd pmos_5p04310591302048_3v1024x8m81_0/S pmos_5p04310591302048_3v1024x8m81_0/S
+ vdd pmos_5p04310591302051_3v1024x8m81_1/S pmos_5p04310591302051_3v1024x8m81_1/S
+ pmos_5p04310591302051_3v1024x8m81
Xnmos_5p04310591302050_3v1024x8m81_0 nmos_5p0431059130208_3v1024x8m81_1/S nmos_5p0431059130208_3v1024x8m81_1/S
+ nmos_5p0431059130208_3v1024x8m81_0/D pmos_5p04310591302051_3v1024x8m81_0/D pmos_5p04310591302051_3v1024x8m81_0/D
+ nmos_5p0431059130208_3v1024x8m81_0/D nmos_5p0431059130208_3v1024x8m81_0/D vss nmos_5p04310591302050_3v1024x8m81
Xnmos_5p04310591302046_3v1024x8m81_0 pmos_5p04310591302051_3v1024x8m81_0/D vss vss
+ vss pmos_5p04310591302051_3v1024x8m81_0/D pmos_5p04310591302051_3v1024x8m81_0/D
+ q pmos_5p04310591302051_3v1024x8m81_0/D q pmos_5p04310591302051_3v1024x8m81_0/D
+ q q pmos_5p04310591302051_3v1024x8m81_0/D vss nmos_5p04310591302046_3v1024x8m81
Xpmos_5p04310591302013_3v1024x8m81_0 nmos_5p0431059130208_3v1024x8m81_1/S nmos_5p0431059130208_3v1024x8m81_1/S
+ se pmos_5p04310591302051_3v1024x8m81_0/D pmos_5p04310591302051_3v1024x8m81_0/D se
+ se vdd pmos_5p04310591302013_3v1024x8m81
Xpmos_5p04310591302049_3v1024x8m81_0 pmos_5p04310591302051_3v1024x8m81_0/D vdd vdd
+ vdd pmos_5p04310591302051_3v1024x8m81_0/D q q pmos_5p04310591302051_3v1024x8m81_0/D
+ q q pmos_5p04310591302051_3v1024x8m81_0/D pmos_5p04310591302051_3v1024x8m81_0/D
+ pmos_5p04310591302051_3v1024x8m81_0/D vdd pmos_5p04310591302049_3v1024x8m81
Xpmos_1p2$$171625516_3v1024x8m81_0 pmos_5p04310591302038_3v1024x8m81_0/D vdd vdd pmos_5p04310591302038_3v1024x8m81_0/D
+ nmos_5p0431059130208_3v1024x8m81_1/S vdd pmos_1p2$$171625516_3v1024x8m81
.ends

.subckt saout_m2_3v1024x8m81 ypass[1] ypass[2] ypass[4] ypass[0] GWEN datain q pcb
+ bb[0] b[0] bb[1] b[2] b[5] b[6] b[7] vss_uq4 vdd vdd_uq2 vdd_uq1 pcb_uq0 pcb_uq1
+ bb[5] mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/bb mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ bb[2] GWE bb[4] WEN bb[7] b[4] men VDD_uq1 VDD b[1] bb[3] ypass[3] ypass[6] ypass[7]
+ VDD_uq0 ypass[5] b[3] vdd_uq3 vdd_uq0 bb[6] vss
Xdin_3v1024x8m81_0 vss datain men sa_3v1024x8m81_0/db sa_3v1024x8m81_0/d sa_3v1024x8m81_0/wep
+ vdd vdd_uq2 pcb_uq0 vss din_3v1024x8m81
Xsacntl_2_3v1024x8m81_0 pcb_uq0 sa_3v1024x8m81_0/se sacntl_2_3v1024x8m81_0/pmos_5p04310591302027_3v1024x8m81_1/S_uq0
+ men sacntl_2_3v1024x8m81_0/pmos_5p04310591302027_3v1024x8m81_2/S_uq0 vdd_uq1 VDD_uq0
+ vss sacntl_2_3v1024x8m81
Xsa_3v1024x8m81_0 sa_3v1024x8m81_0/qp sa_3v1024x8m81_0/qn sa_3v1024x8m81_0/wep sa_3v1024x8m81_0/se
+ pcb_uq0 sa_3v1024x8m81_0/db vdd_uq2 vdd sa_3v1024x8m81_0/d vss sa_3v1024x8m81
Xmux821_3v1024x8m81_0 b[6] bb[6] bb[5] sa_3v1024x8m81_0/db sa_3v1024x8m81_0/d sa_3v1024x8m81_0/db
+ ypass[0] b[1] ypass[1] ypass[3] mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/bb
+ bb[4] ypass[5] sa_3v1024x8m81_0/d b[5] bb[3] ypass[2] ypass[4] b[4] ypass[6] sa_3v1024x8m81_0/d
+ ypass[7] b[7] sa_3v1024x8m81_0/d bb[7] sa_3v1024x8m81_0/d bb[2] bb[1] sa_3v1024x8m81_0/db
+ sa_3v1024x8m81_0/db sa_3v1024x8m81_0/d ypass[3] ypass[7] ypass[2] ypass[0] b[3]
+ vdd_uq0 ypass[5] ypass[1] ypass[4] sa_3v1024x8m81_0/d mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ b[2] vdd_uq3 vss ypass[6] sa_3v1024x8m81_0/d pcb_uq0 mux821_3v1024x8m81
Xwen_wm1_3v1024x8m81_0 GWEN men sa_3v1024x8m81_0/wep VDD_uq1 WEN vss VDD wen_wm1_3v1024x8m81
Xoutbuf_oe_3v1024x8m81_0 sa_3v1024x8m81_0/qp sa_3v1024x8m81_0/qn sa_3v1024x8m81_0/se
+ q GWE vss vdd outbuf_oe_3v1024x8m81
.ends

.subckt x018SRAM_cell1_3v1024x8m81 m3_82_330# a_248_342# a_248_592# a_62_178# w_30_512#
+ a_430_96# a_110_96# VSUBS
X0 a_248_592# a_192_298# a_110_250# w_30_512# pfet_03v3 ad=0.1613p pd=1.39u as=0.1238p ps=1.44u w=0.28u l=0.28u
X1 a_248_342# a_192_298# a_110_250# VSUBS nfet_03v3 ad=0.171p pd=1.33u as=0.15665p ps=1.32u w=0.45u l=0.28u
X2 a_192_298# a_110_250# a_248_592# w_30_512# pfet_03v3 ad=0.1238p pd=1.44u as=0.1613p ps=1.39u w=0.28u l=0.28u
X3 a_192_298# a_110_250# a_248_342# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.171p ps=1.33u w=0.45u l=0.28u
X4 a_110_250# a_62_178# a_110_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
X5 a_192_298# a_62_178# a_430_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
.ends

.subckt x018SRAM_cell1_2x_3v1024x8m81 018SRAM_cell1_3v1024x8m81_0/a_62_178# 018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_62_178# 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_3v1024x8m81_1/a_248_342# VSUBS
X018SRAM_cell1_3v1024x8m81_1 018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_3v1024x8m81_1/a_248_592# 018SRAM_cell1_3v1024x8m81_1/a_62_178# 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_3v1024x8m81_1/a_110_96# VSUBS
+ x018SRAM_cell1_3v1024x8m81
X018SRAM_cell1_3v1024x8m81_0 018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_3v1024x8m81_0/a_62_178# 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_3v1024x8m81_1/a_110_96# VSUBS
+ x018SRAM_cell1_3v1024x8m81
.ends

.subckt rarray4_1024_3v1024x8m81 m3_n1397_74227# m3_n1397_30097# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ m3_n1397_64531# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ m3_n1397_39793# m3_n1397_41503# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ m3_n1397_48775# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2221# m3_n1397_61609# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ m3_n1397_70591# m3_n1397_26461# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# m3_n1397_53125#
+ m3_n1397_17977# m3_n1397_51913# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ m3_n1397_8779# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# m3_n1397_31309# m3_n1397_76153# m3_n1397_40291# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ m3_n1397_49987# m3_n1397_16765# m3_n1397_3433# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# m3_n1397_20401# m3_n1397_1009# m3_n1397_70093# m3_n1397_57259# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ m3_n1397_62107# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# m3_n1397_54337#
+ m3_n1397_19687# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# m3_n1397_71305# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96# m3_n1397_60895#
+ m3_n1397_48277# m3_n1397_36655# m3_n1397_59185# m3_n1397_9991# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# m3_n1397_27673#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ m3_n1397_57973# m3_n1397_68881# m3_n1397_13129# m3_n1397_51199# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74941# m3_n1397_35443# m3_n1397_20899# m3_n1397_43429# m3_n1397_53623#
+ m3_n1397_12415# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# m3_n1397_41005#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96# m3_n1397_73729#
+ m3_n1397_23323# m3_n1397_77365# m3_n1397_52411# m3_n1397_37369# m3_n1397_14839#
+ m3_n1397_15553# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11917# m3_n1397_5857# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ m3_n1397_34231# m3_n1397_69379# m3_n1397_14341# m3_n1397_19189# m3_n1397_10705#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96# m3_n1397_4645#
+ m3_n1397_67669# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22825# m3_n1397_68167# m3_n1397_38581# m3_n1397_36157# m3_n1397_56047#
+ m3_n1397_21613# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ m3_n1397_73015# m3_n1397_247# m3_n1397_56761# m3_n1397_28171# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# m3_n1397_1507# m3_n1397_63319# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# m3_n1397_47065#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# m3_n1397_24037#
+ m3_n1397_64033# m3_n1397_29383# m3_n1397_46351# m3_n1397_34945# m3_n1397_72517#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# m3_n1397_37867#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# m3_n1397_50701#
+ m3_n1397_9493# m3_n1397_54835# m3_n1397_8281# m3_n1397_17263# m3_n1397_31807# m3_n1397_65743#
+ m3_n1397_71803# m3_n1397_76651# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49489# m3_n1397_5143# m3_n1397_55549# m3_n1397_28885# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# m3_n1397_33019# m3_n1397_45853# m3_n1397_62821# m3_n1397_33733# m3_n1397_42715#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ m3_n1397_44641# m3_n1397_58471# m3_n1397_45139# m3_n1397_7069# m3_n1397_39079# m3_n1397_30595#
+ m3_n1397_7567# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ m3_n1397_16051# m3_n1397_25249# m3_n1397_65245# m3_n1397_3931# m3_n1397_42217# m3_n1397_43927#
+ m3_n1397_75439# m3_n1397_25747# m3_n1397_11203# m3_n1397_66457# m3_n1397_24535#
+ m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ VSUBS m3_n1397_60397#
X018SRAM_cell1_2x_3v1024x8m81_362 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_395 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_351 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_340 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_384 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_373 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1417 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1406 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1439 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1428 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_192 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_181 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_170 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1984 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1962 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1951 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1973 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1940 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1995 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1258 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1225 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1214 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1247 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1269 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1236 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1203 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1792 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_906 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_917 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1770 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1781 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_928 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_939 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1011 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1000 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1088 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1066 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1033 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1055 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1077 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1044 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1022 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1099 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_725 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_758 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_736 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_747 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_714 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_703 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_769 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_588 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_544 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_533 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_555 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_599 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_566 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_577 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_500 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_511 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_522 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_363 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_330 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_341 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_396 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_352 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_374 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_385 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1418 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1407 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1429 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_193 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_182 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_160 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_171 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1952 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1985 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1930 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1974 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1941 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1996 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1963 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1204 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1248 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1226 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1215 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1237 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1259 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1760 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1793 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_907 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_918 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_929 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1782 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1771 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1034 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1001 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1045 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1023 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1012 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1056 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1089 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1078 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1067 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1590 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_737 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_759 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_748 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_726 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_715 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_704 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_512 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_589 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_578 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_534 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_556 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_545 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_567 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_523 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_501 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_320 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_342 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_331 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_364 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_386 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_397 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_353 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_375 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1408 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1419 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_183 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_161 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_172 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_150 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_194 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1920 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1942 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1931 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1986 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1953 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1975 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1997 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1964 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1216 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1205 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1227 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1249 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1238 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1761 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1783 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1750 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1772 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1794 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_919 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_908 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1057 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1002 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1079 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1046 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1024 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1035 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1068 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1013 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1591 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1580 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_727 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_749 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_738 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_716 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_705 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_524 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_513 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_502 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_579 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_535 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_546 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_557 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_568 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_365 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_354 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_310 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_376 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_343 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_321 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_332 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_387 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_398 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1409 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_184 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_195 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_162 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_173 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_151 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_140 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1954 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1921 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1976 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1943 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1910 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1965 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1932 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1987 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1998 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1217 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1239 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1206 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1228 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1762 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1795 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1784 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1751 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1773 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1740 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_909 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1058 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1025 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1003 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1047 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1069 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1036 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1014 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1570 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1592 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_706 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1581 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_728 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_739 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_717 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_547 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_536 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_558 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_525 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_514 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_503 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_569 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_388 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_333 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_300 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_399 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_344 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_311 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_377 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_366 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_322 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_355 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_196 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_185 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_163 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_174 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_152 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_141 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_130 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1922 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1988 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1955 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1944 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1977 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1911 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1999 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1966 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1933 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1900 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1218 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1207 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1229 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1730 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1796 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1763 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1752 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1785 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1774 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1741 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1026 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1059 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1004 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1048 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1037 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1015 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1571 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_729 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_718 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1560 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1593 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_707 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1582 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1390 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_548 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_537 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_559 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_526 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_515 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_504 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_389 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_334 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_301 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_345 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_378 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_367 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_323 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_312 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_356 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_890 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_120 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_131 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_197 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_186 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_164 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_175 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_153 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_142 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1956 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1923 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1989 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1978 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1912 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1945 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1934 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1967 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1901 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1219 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1208 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1731 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1720 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1764 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1797 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1786 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1753 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1742 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1775 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1027 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1005 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1016 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1049 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1038 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1572 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1561 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1550 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1583 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_719 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1594 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_708 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1380 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1391 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_549 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_538 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_527 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_516 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_505 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_302 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_324 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_313 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_335 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_379 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_346 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_368 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_357 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_880 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_891 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_165 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_143 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_121 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_110 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_154 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_132 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_198 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_187 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_176 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1924 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1913 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1902 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1957 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1946 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1979 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1968 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1935 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1209 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1732 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1765 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1754 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1721 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1710 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1743 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1798 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1787 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1776 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1028 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1006 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1039 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1017 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1540 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1573 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1562 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1595 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1584 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1551 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_709 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1381 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1370 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_506 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1392 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_539 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_528 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_517 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_303 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_347 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_336 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_325 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_314 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_358 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_369 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_892 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_881 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_870 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_188 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_199 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_166 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_177 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_144 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_111 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_100 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_133 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_122 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_155 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1958 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1925 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1914 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1947 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1936 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1903 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1969 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1700 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1766 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1733 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1799 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1788 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1722 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1755 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1777 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1744 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1711 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1029 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1007 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1018 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1574 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1541 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1596 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1530 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1563 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1585 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1552 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1382 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_529 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1371 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_507 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_518 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1393 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1360 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1190 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_304 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_348 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_326 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_337 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_315 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_359 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_893 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_882 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_871 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_860 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_167 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_189 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_178 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_112 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_134 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_156 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_145 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_101 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_123 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1926 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1959 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1948 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1915 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1937 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1904 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_690 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1734 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1701 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1767 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1756 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1789 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1723 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1778 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1745 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1712 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1019 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1008 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1531 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1520 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1542 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1575 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1564 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1597 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1586 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1553 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1350 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1383 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1372 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2040 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1361 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_508 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_519 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1394 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1191 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1180 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_305 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_327 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_349 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_338 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_316 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_894 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_872 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_883 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_850 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_861 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_113 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_102 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_168 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_179 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_135 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_157 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_146 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_124 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1927 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1916 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1949 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1938 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1905 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_691 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_680 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1702 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1713 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1735 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1768 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1724 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1757 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1746 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1779 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1009 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1510 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1543 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1532 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1565 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1554 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1521 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1576 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1598 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1587 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1351 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1384 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1340 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1373 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2041 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1362 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1395 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2030 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_509 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1192 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_306 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1181 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1170 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_328 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_339 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_317 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_840 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_851 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_862 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_895 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_873 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_884 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_114 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_136 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_147 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_103 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_125 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_169 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_158 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1906 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1928 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1917 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1939 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_692 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_681 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_670 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1703 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1736 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1725 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1714 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1747 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1769 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1758 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1511 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1544 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1577 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1500 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1566 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1599 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1533 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1588 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1522 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1555 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2020 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2042 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2031 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1352 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1385 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1374 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1341 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1396 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1363 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1330 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1160 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1193 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_329 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1182 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_307 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_318 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1171 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_874 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_885 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_830 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_841 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_852 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_863 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_896 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_115 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_159 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_148 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_104 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_126 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_137 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1929 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1918 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1907 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_693 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_682 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_660 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_671 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1704 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1737 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1726 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1759 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1748 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1715 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_490 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1512 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1578 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1545 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1534 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1567 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1501 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1589 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1556 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1523 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2021 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1320 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2010 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2043 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1331 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2032 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1386 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1353 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1342 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1375 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1397 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1364 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1161 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1150 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1172 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1194 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_319 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1183 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_308 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_897 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_875 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_886 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_831 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_842 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_853 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_820 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_864 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_116 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_127 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_149 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_105 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_138 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1919 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1908 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_694 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_650 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_683 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_661 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_672 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1738 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1705 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1727 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1749 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1716 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_480 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_491 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1513 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1502 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1568 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1546 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1535 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1557 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1524 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1579 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2022 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1321 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1354 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2044 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1310 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1343 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2011 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1365 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1332 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2033 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2000 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1376 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1398 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1387 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1184 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1162 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1151 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1173 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1140 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1195 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_309 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_810 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_898 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_876 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_887 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_843 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_832 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_854 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_821 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_865 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_106 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_128 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_117 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_139 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1909 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_651 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_640 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_695 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_662 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_684 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_673 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1728 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1706 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1717 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1739 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_470 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_481 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_492 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1536 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1514 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1503 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1525 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1547 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1569 m3_n1397_59683# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_59683# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_60397#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1558 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1344 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1377 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2023 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1322 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2012 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1311 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2045 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1366 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1333 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1300 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2034 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2001 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1388 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1355 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1399 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1152 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1185 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1130 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1174 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1141 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1196 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1163 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_833 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_844 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_800 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_811 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_822 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_899 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_877 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_888 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_855 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_866 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_118 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_107 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_129 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_630 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_652 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_641 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_663 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_685 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_674 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_696 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1729 m3_n1397_65743# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_65743# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_66457#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1718 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1707 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_471 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_460 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_482 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_493 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1504 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1537 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1559 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1526 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1548 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1515 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_290 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2024 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_90 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2013 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2002 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1378 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1312 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1345 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2046 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1367 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1334 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1301 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2035 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1389 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1356 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1323 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1890 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1120 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1131 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1186 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1153 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1175 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1142 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1197 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1164 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_834 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_801 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_845 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_856 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_867 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_812 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_823 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_878 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_889 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_108 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_119 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_631 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_620 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_653 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_642 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_686 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_697 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_675 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_664 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1719 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1708 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_472 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_461 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_450 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_494 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_483 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1538 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1505 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1527 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1549 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1516 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_280 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_291 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_91 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_80 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1313 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2025 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2014 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2047 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1302 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2036 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2003 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1346 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1379 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1368 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1335 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1357 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1324 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1891 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1880 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1154 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1121 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1143 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1110 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1132 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1187 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1176 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1198 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1165 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_879 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_835 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_824 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_802 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_813 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_846 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_868 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_857 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_109 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_621 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_610 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_654 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_643 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_687 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_632 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_698 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_676 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_665 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1709 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_451 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_440 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_495 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_484 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_462 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_473 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_4 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1506 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1539 m3_n1397_58471# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_58471# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_59185#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1528 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1517 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_292 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_281 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_270 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_92 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_70 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_81 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1314 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1347 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2026 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2015 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1336 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1303 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2037 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2004 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1325 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1369 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1358 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1892 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1881 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1870 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1122 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1188 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1155 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1144 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1177 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1111 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1166 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1133 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1100 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1199 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_825 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_803 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_814 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_836 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_847 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_858 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_869 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_622 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_611 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_600 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_633 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_688 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_644 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_677 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_699 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_666 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_655 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_452 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_430 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_463 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_441 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_485 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_474 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_496 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_5 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1507 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1529 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1518 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_260 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_282 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_293 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_271 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_93 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_60 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_82 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_71 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2016 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1348 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1315 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1304 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1337 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2038 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2005 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1359 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1326 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2027 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1860 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1893 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1882 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1871 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1156 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1123 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1189 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1178 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1112 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1145 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1134 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1167 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1101 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1690 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_826 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_804 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_815 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_837 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_859 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_848 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_623 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_612 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_601 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_634 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_667 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_645 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_656 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_689 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_678 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_464 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_475 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_453 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_497 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_420 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_431 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_442 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_486 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_6 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1508 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1519 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_261 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_283 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_250 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_294 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_272 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_50 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_94 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2006 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_61 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_72 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_83 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2017 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1316 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1349 m3_n1397_51199# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_51199# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_51913#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1338 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1305 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2039 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1327 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2028 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1894 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1861 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1850 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1883 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1872 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1113 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1102 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1124 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1157 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1146 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1179 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1168 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1135 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1691 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1680 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_816 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_838 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_827 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_805 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_849 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_624 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_602 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_613 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_635 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_679 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_657 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_668 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_646 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_476 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_454 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_421 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_498 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_465 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_410 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_443 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_432 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_487 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_7 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1509 m3_n1397_57259# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_57259# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_57973#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_251 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_240 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_262 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_284 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_295 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_273 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_40 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_51 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_62 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_73 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_84 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2018 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_95 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2007 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2029 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1317 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1306 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1339 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1328 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1851 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1840 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1862 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1895 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1884 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1873 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1125 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1114 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1136 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1103 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1158 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1147 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1169 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1670 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1692 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1681 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_817 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_839 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_828 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_806 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_625 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_603 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_614 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_636 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_658 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_669 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_647 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_422 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_411 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_433 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_400 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_477 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_455 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_499 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_466 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_444 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_488 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_8 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_230 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_263 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_252 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_241 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_274 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_296 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_285 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_41 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_52 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_30 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_96 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_63 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_74 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_85 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2019 m3_n1397_76651# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_76651# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_77365#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1318 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1307 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2008 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1329 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1830 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1863 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1852 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1874 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1841 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1896 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1885 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1126 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1159 m3_n1397_43927# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_43927# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_44641#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1148 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1115 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1137 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1104 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1671 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1660 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1693 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1682 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_818 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_829 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_807 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_604 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_615 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1490 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_626 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_648 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_659 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_637 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_467 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_456 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_423 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_412 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_434 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_445 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_401 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_478 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_489 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_9 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_990 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_220 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_231 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_297 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_286 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_253 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_275 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_242 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_264 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_42 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_53 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_20 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_31 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_64 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_75 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_86 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_97 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1319 m3_n1397_49987# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_49987# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_50701#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1308 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2009 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1831 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1864 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1897 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1820 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1886 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1853 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1842 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1875 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1127 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1116 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1149 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1138 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1105 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1672 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1694 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1661 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1683 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1650 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_808 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_819 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1480 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_627 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_605 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_616 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_649 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_638 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1491 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_457 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_424 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_413 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_468 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_435 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_446 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_479 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_402 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_980 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_991 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_221 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_210 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_298 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_287 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_254 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_276 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_243 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_265 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_232 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_10 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_21 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_32 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_43 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_54 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_65 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_87 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_98 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_76 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1309 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1832 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1898 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1865 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1854 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1887 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1821 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1876 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1810 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1843 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1128 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1117 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1106 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1139 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1640 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1673 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1662 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1695 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1684 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1651 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_809 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1481 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1470 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1492 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_628 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_606 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_617 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_639 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_425 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_414 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_469 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_447 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_458 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_436 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_403 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_981 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_992 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_970 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_200 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_222 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_211 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_233 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_299 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_288 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_255 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_277 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_244 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_266 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_44 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_11 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_55 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_22 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_33 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_66 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_99 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_88 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_77 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1800 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1833 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1822 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1811 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1888 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1866 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1855 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1877 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1844 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1899 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1118 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1107 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1129 m3_n1397_42715# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_42715# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_43429#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1641 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1674 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1630 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1663 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1652 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1696 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1685 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1482 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1471 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1493 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1460 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_607 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_629 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_618 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1290 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_415 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_404 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_448 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_426 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_437 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_459 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_960 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_971 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_982 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_993 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_201 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_234 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_223 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_256 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_245 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_212 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_278 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_289 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_267 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_790 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_45 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_12 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_34 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_23 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_56 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_67 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_78 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_89 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1856 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1834 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1801 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1823 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1845 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1812 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1889 m3_n1397_71803# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_71803# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_72517#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1878 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1867 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1119 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1108 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1664 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1697 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1642 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1631 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1686 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1653 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1620 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1675 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1472 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1450 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1494 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1461 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1483 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_608 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_619 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1280 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_449 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_416 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_438 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_405 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_427 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1291 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_983 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_961 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_950 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_994 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_972 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_235 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_202 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_257 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_279 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_246 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_268 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_224 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_213 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_791 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_780 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_46 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_13 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_35 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_24 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_57 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_68 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_79 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1824 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1857 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1802 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1879 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1846 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1813 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1868 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1835 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1109 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1698 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1632 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1665 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1610 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1687 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1654 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1621 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1676 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1643 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1440 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1473 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_609 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1495 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1462 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1484 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1451 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1281 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1270 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1292 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_439 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_417 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_406 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_428 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_940 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_984 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_962 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_951 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_995 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_973 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_203 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_258 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_269 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_247 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_214 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_225 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_236 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_781 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_792 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_770 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_14 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_47 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_36 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_25 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_58 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_69 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1858 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1825 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1847 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1814 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1869 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1836 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1803 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1600 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1622 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1611 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1666 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1633 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1699 m3_n1397_64531# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_64531# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_65245#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1688 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1655 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1677 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1644 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1474 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1441 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1463 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1430 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1452 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1496 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1485 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1282 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1271 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1293 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1260 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_418 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_429 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_407 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_941 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_985 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_930 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_963 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_996 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_974 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_952 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1090 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_204 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_215 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_226 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_259 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_248 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_237 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_760 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_782 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_793 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_771 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_15 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_48 m3_n1397_6355# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_7069#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_37 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_26 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_59 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1815 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1804 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1826 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1859 m3_n1397_70591# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_70591# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_71305#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1848 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1837 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_590 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1634 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1601 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1656 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1623 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1645 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1612 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1667 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1689 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1678 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1442 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1475 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1464 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1497 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1431 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1486 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1453 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1420 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1250 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1283 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1272 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1294 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1261 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_419 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_408 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_920 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_942 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_931 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_953 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_986 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_997 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_964 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_975 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_975/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_216 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1091 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_205 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_227 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_238 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1080 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_249 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_761 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_750 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_783 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_794 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_772 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_49 m3_n1397_7567# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_8281#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_38 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_27 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_16 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1827 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1816 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1838 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1805 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1849 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_591 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_580 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1602 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1668 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1635 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1624 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1657 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1679 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1646 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1613 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1410 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1476 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1443 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1498 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1432 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1465 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1454 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1487 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1421 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1240 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1284 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1251 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1273 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_409 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1262 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1295 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_921 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_910 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_943 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_965 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_976 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_932 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_954 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_987 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_998 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1081 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1070 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_217 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1092 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_206 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_239 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_228 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_762 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_751 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_740 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_784 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_773 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_98/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_795 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_39 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_17 m3_n1397_1507# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_2221#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_28 m3_n1397_3931# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_4645#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1828 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1817 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1806 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1839 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_592 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_581 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_570 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1636 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1603 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1669 m3_n1397_63319# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_63319# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_64033#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1658 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1625 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1614 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1647 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1411 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1400 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1422 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1444 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1477 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1466 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1499 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1433 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1488 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1455 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1252 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1241 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1230 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1263 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1285 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1274 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1296 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_900 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_922 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_944 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_988 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_911 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_999 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_966 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_977 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_933 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_955 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1060 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1093 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1082 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1071 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_207 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_218 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_229 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_763 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_752 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_730 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_741 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_785 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_774 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_796 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_18 m3_n1397_247# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_1009#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_29 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1829 m3_n1397_69379# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_69379# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_70093#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1818 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1807 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_560 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_593 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_582 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_571 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1604 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1637 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1626 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1659 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1648 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1615 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_390 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1412 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1445 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1434 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1401 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1456 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1423 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1478 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1467 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1489 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1990 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1220 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1286 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1253 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1242 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1275 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1297 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1264 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1231 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_901 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_934 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_923 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_945 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_989 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_912 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_967 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_967/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_978 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_956 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1094 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1061 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1050 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1083 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1072 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_208 m3_n1397_8779# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_9493#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_219 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_731 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_742 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_720 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_764 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_753 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_786 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_775 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_797 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_19 m3_n1397_2719# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_3433#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1819 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1808 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_550 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_583 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_561 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_572 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_594 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1638 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1605 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1627 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1616 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1649 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_391 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_380 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1446 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1413 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1479 m3_n1397_56047# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_56047# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_56761#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1468 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1402 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1435 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1457 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1424 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1991 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1980 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1254 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1221 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1287 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1276 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1210 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1243 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1298 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1265 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1232 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_902 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_935 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_924 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_913 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_946 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_968 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_979 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_957 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1062 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_209 m3_n1397_9991# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_10705#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1095 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1084 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1051 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1040 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1073 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_765 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_743 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_721 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_754 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_732 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_710 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_776 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_787 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_798 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1809 m3_n1397_68167# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_68167# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_68881#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_551 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_540 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_584 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_562 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_573 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_595 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1606 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1639 m3_n1397_62107# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_62107# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_62821#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1628 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1617 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_392 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_370 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_381 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1414 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1447 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1436 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1469 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1403 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1458 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1425 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1992 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1981 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1970 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1222 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1211 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1200 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1255 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1288 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1244 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1277 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1266 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1299 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1233 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_903 m3_n1397_36655# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_36655# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_37369#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_936 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_925 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_947 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_914 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_958 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_969 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1030 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1063 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1052 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1041 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_977/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1096 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1085 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1074 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_766 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_744 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_755 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_733 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_722 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_700 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_711 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_999/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_788 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_777 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_799 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_541 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_530 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_552 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_563 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_585 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_574 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_596 m3_n1397_33019# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_33019# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_33733#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1607 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1629 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1618 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_360 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_371 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_393 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_382 m3_n1397_13627# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_14341#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1404 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1415 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1448 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1437 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1426 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1459 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_190 m3_n1397_11203# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_11917#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1960 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1993 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1982 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1971 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1223 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1212 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1245 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1234 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1201 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_979/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1256 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1289 m3_n1397_48775# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_48775# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_49489#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1278 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1267 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1790 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_904 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_937 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_926 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_915 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_959 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_99/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_948 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1031 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1064 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1097 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1086 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1053 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1042 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1075 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1020 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_701 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_745 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_767 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_756 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_734 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_723 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_712 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_778 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_789 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_542 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_531 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_520 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_553 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_586 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_564 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_575 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_597 m3_n1397_34231# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_34231# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_34945#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1608 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1619 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_361 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_394 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_350 m3_n1397_5143# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_5857#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_372 m3_n1397_17263# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_17977#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_383 m3_n1397_14839# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_15553#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1416 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1438 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1405 m3_n1397_52411# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_52411# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_53125#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1427 m3_n1397_53623# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_53623# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_54337#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1449 m3_n1397_54835# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_54835# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_55549#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_191 m3_n1397_12415# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_13129#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_180 m3_n1397_16051# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_16765#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1961 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1994 m3_n1397_75439# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_75439# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_76153#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1950 m3_n1397_73015# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_73015# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_73729#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1983 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1972 m3_n1397_74227# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_74227# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_74941#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1224 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1257 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1246 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1279 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1213 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1268 m3_n1397_47563# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_47563# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_48277#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1202 m3_n1397_45139# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_45139# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_45853#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1235 m3_n1397_46351# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_971/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_46351# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_47065#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1791 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1780 m3_n1397_66955# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_66955# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_67669#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_927 m3_n1397_31807# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_31807# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_32521#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_905 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_916 m3_n1397_35443# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_35443# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_36157#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_938 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_65/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_949 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1032 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1010 m3_n1397_18475# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_96/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_19189#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1098 m3_n1397_41503# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_81/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_41503# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_42217#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1065 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1054 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_719/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1087 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_717/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1076 m3_n1397_40291# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_40291# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_41005#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1043 m3_n1397_39079# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_39079# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_39793#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1021 m3_n1397_19687# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_19687# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_20401#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_724 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_713 m3_n1397_29383# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_713/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_29383# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_30097#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_702 m3_n1397_28171# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_973/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_28171# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_28885#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_746 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_757 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_735 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_779 m3_n1397_26959# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_82/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_26959# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_27673#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_768 m3_n1397_24535# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_24535# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_25249#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_543 m3_n1397_25747# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_25747# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_26461#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_532 m3_n1397_22111# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_993/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_22111# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_22825#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_565 m3_n1397_23323# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_23323# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_24037#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_576 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_554 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_997/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_521 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_965/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_510 m3_n1397_20899# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_969/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_20899# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_21613#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_587 m3_n1397_30595# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_995/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_30595# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_31309#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_598 m3_n1397_37867# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_715/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_37867# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_38581#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1609 m3_n1397_60895# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609# 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_2x_3v1024x8m81_89/018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ m3_n1397_60895# VSUBS 018SRAM_strap1_bndry_3v1024x8m81_9/w_91_512# m3_n1397_61609#
+ VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
.ends

.subckt dcap_103_novia_3v1024x8m81 w_n205_0# a_n30_42# a_n119_86#
X0 a_n119_86# a_n30_42# a_n119_86# w_n205_0# pfet_03v3 ad=0.4717p pd=3.01u as=0 ps=0 w=1.06u l=1.74u
.ends

.subckt pmos_5p04310591302095_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.4251p pd=2.155u as=0.7194p ps=4.15u w=1.635u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.7194p pd=4.15u as=0.4251p ps=2.155u w=1.635u l=0.28u
.ends

.subckt x018SRAM_cell1_dummy_R_3v1024x8m81 m3_82_330# a_248_342# a_62_178# w_30_512#
+ a_430_96# a_110_96# a_192_298# VSUBS
X0 a_192_298# a_192_298# a_110_250# w_30_512# pfet_03v3 ad=0.1613p pd=1.39u as=0.1238p ps=1.44u w=0.28u l=0.28u
X1 a_248_342# a_192_298# a_110_250# VSUBS nfet_03v3 ad=0.171p pd=1.33u as=0.15665p ps=1.32u w=0.45u l=0.28u
X2 a_408_342# a_248_342# a_192_298# w_30_512# pfet_03v3 ad=0.1238p pd=1.44u as=0.1613p ps=1.39u w=0.28u l=0.28u
X3 a_408_342# a_248_342# a_248_342# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.171p ps=1.33u w=0.45u l=0.28u
X4 a_110_250# a_62_178# a_110_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
X5 a_408_342# a_62_178# a_430_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
.ends

.subckt x018SRAM_cell1_dummy_3v1024x8m81 m3_82_330# a_248_342# a_248_592# w_82_512#
+ a_62_178# m2_346_89# m2_134_89# VSUBS
X0 a_248_592# a_192_298# a_110_250# w_82_512# pfet_03v3 ad=0.1613p pd=1.39u as=0.1238p ps=1.44u w=0.28u l=0.28u
X1 a_248_342# a_192_298# a_110_250# VSUBS nfet_03v3 ad=0.171p pd=1.33u as=0.15665p ps=1.32u w=0.45u l=0.28u
X2 a_192_298# a_110_250# a_248_592# w_82_512# pfet_03v3 ad=0.1238p pd=1.44u as=0.1613p ps=1.39u w=0.28u l=0.28u
X3 a_192_298# a_110_250# a_248_342# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.171p ps=1.33u w=0.45u l=0.28u
X4 a_110_250# a_62_178# a_110_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
X5 a_192_298# a_62_178# a_430_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
.ends

.subckt pmos_5p04310591302097_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=1.2909p pd=5.485u as=2.1846p ps=10.81u w=4.965u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=2.1846p pd=10.81u as=1.2909p ps=5.485u w=4.965u l=0.28u
.ends

.subckt nmos_5p04310591302096_3v1024x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=1.0309p pd=4.485u as=1.7446p ps=8.81u w=3.965u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=1.7446p pd=8.81u as=1.0309p ps=4.485u w=3.965u l=0.28u
.ends

.subckt ypass_gate_3v1024x8m81_0 vss bb db ypass d pcb vdd_uq0 m3_0_2091# pmos_5p0431059130201_3v1024x8m81_2/D
+ m3_0_2831# a_64_1295# m3_0_3056# pmos_5p0431059130201_3v1024x8m81_0/D m3_0_3781#
+ m3_0_1632# VSUBS m3_0_3536# b m3_0_3291# m3_0_2331# vdd m3_0_2581#
Xnmos_5p0431059130200_3v1024x8m81_0 pmos_5p0431059130201_3v1024x8m81_2/D a_64_1295#
+ bb VSUBS nmos_5p0431059130200_3v1024x8m81
Xnmos_5p0431059130200_3v1024x8m81_1 pmos_5p0431059130201_3v1024x8m81_0/D a_64_1295#
+ b VSUBS nmos_5p0431059130200_3v1024x8m81
Xpmos_5p0431059130201_3v1024x8m81_0 pmos_5p0431059130201_3v1024x8m81_0/D nmos_5p0431059130202_3v1024x8m81_0/D
+ vdd_uq0 b pmos_5p0431059130201_3v1024x8m81
Xpmos_5p0431059130201_3v1024x8m81_1 b pcb vdd bb pmos_5p0431059130201_3v1024x8m81
Xpmos_5p0431059130201_3v1024x8m81_2 pmos_5p0431059130201_3v1024x8m81_2/D nmos_5p0431059130202_3v1024x8m81_0/D
+ vdd bb pmos_5p0431059130201_3v1024x8m81
Xnmos_5p0431059130202_3v1024x8m81_0 nmos_5p0431059130202_3v1024x8m81_0/D a_64_1295#
+ a_64_1295# VSUBS VSUBS VSUBS nmos_5p0431059130202_3v1024x8m81
X0 vdd pcb b vdd pfet_03v3 ad=0.94105p pd=4.37u as=0.51437p ps=2.24u w=1.595u l=0.28u
X1 bb pcb vdd vdd pfet_03v3 ad=0.51437p pd=2.24u as=1.13245p ps=4.61u w=1.595u l=0.28u
X2 nmos_5p0431059130202_3v1024x8m81_0/D a_64_1295# vdd_uq0 vdd_uq0 pfet_03v3 ad=0.1946p pd=1.255u as=0.38225p ps=2.49u w=0.695u l=0.28u
X3 vdd_uq0 a_64_1295# nmos_5p0431059130202_3v1024x8m81_0/D vdd_uq0 pfet_03v3 ad=0.50735p pd=2.85u as=0.1946p ps=1.255u w=0.695u l=0.28u
X4 b pcb vdd vdd pfet_03v3 ad=0.51437p pd=2.24u as=1.13245p ps=4.61u w=1.595u l=0.28u
X5 vdd pcb bb vdd pfet_03v3 ad=0.94105p pd=4.37u as=0.51437p ps=2.24u w=1.595u l=0.28u
.ends

.subckt nmos_5p04310591302098_3v1024x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.1664p pd=1.16u as=0.2816p ps=2.16u w=0.64u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.2816p pd=2.16u as=0.1664p ps=1.16u w=0.64u l=0.28u
.ends

.subckt rdummy_3v512x4_3v1024x8m81 018SRAM_cell1_dummy_R_3v1024x8m81_63/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v1024x8m81_57/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_24/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_42/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_30/m2_346_89# 018SRAM_cell1_2x_3v1024x8m81_42/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_129/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_13/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_58/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_dummy_3v1024x8m81_30/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_113/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_13/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_129/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_58/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_121/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_34/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_73/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_73/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_34/a_248_342# 018SRAM_cell1_dummy_3v1024x8m81_40/m2_346_89#
+ pmos_5p04310591302097_3v1024x8m81_0/D 018SRAM_cell1_2x_3v1024x8m81_45/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_37/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_11/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_63/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ m3_15667_n5798# 018SRAM_cell1_dummy_3v1024x8m81_40/m2_134_89# 018SRAM_cell1_2x_3v1024x8m81_11/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_43/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_83/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_44/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_43/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_59/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_83/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_44/a_248_342# 018SRAM_cell1_dummy_3v1024x8m81_50/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_11/m2_346_89# 018SRAM_cell1_2x_3v1024x8m81_59/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_2/m2_346_89# 018SRAM_cell1_2x_3v1024x8m81_13/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_dummy_3v1024x8m81_50/m2_134_89# 018SRAM_cell1_2x_3v1024x8m81_36/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_3v1024x8m81_2/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_11/m2_134_89#
+ 018SRAM_cell1_2x_3v1024x8m81_41/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_41/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_1/a_248_592# 018SRAM_cell1_dummy_R_3v1024x8m81_38/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_93/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_54/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_57/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_12/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_15/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_93/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_54/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_57/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_12/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v1024x8m81_60/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_15/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_57/a_192_298#
+ 018SRAM_cell1_dummy_3v1024x8m81_21/m2_346_89# 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_3/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_60/m2_134_89# 018SRAM_cell1_dummy_R_3v1024x8m81_127/w_30_512#
+ 018SRAM_cell1_dummy_3v1024x8m81_21/m2_134_89# w_15880_n13729# 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_9/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_44/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_9/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_10/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_64/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_25/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_10/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_34/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_60/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v1024x8m81_67/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_25/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_3/018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_64/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_31/m2_346_89# 018SRAM_cell1_dummy_R_3v1024x8m81_67/a_192_298#
+ 018SRAM_cell1_2x_3v1024x8m81_42/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_42/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_58/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_31/m2_134_89# 018SRAM_cell1_dummy_R_3v1024x8m81_123/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_58/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_74/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_25/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_35/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v1024x8m81_74/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_40/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_35/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_77/a_192_298# 018SRAM_cell1_dummy_3v1024x8m81_41/m2_346_89#
+ 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_1/a_248_592# 018SRAM_cell1_2x_3v1024x8m81_40/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_38/a_192_298#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_63/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_56/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_41/m2_134_89# 018SRAM_cell1_2x_3v1024x8m81_11/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_11/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_56/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_84/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_45/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_84/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_45/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_12/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_3v1024x8m81_3/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_51/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_87/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_43/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_3v1024x8m81_12/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_3/m2_134_89#
+ 018SRAM_cell1_2x_3v1024x8m81_59/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v1024x8m81_100/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_51/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_12/m2_134_89#
+ 018SRAM_cell1_2x_3v1024x8m81_41/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_25/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_100/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_4/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_94/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_25/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_103/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_41/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_55/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_57/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_94/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_16/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_57/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_55/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_16/a_248_342# 018SRAM_cell1_dummy_3v1024x8m81_61/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_22/m2_346_89# 018SRAM_cell1_dummy_R_3v1024x8m81_97/a_192_298#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_58/a_192_298# ypass_gate_3v1024x8m81_0_0/vss 018SRAM_cell1_2x_3v1024x8m81_11/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_dummy_3v1024x8m81_61/m2_134_89# 018SRAM_cell1_dummy_R_3v1024x8m81_110/m3_82_330#
+ m1_16100_n16182# 018SRAM_cell1_dummy_3v1024x8m81_22/m2_134_89# 018SRAM_cell1_2x_3v1024x8m81_48/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_110/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_113/a_192_298#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_65/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_10/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_26/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_10/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_65/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_77/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_26/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_32/m2_346_89# 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_120/m3_82_330# 018SRAM_cell1_dummy_3v1024x8m81_32/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_120/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_42/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_123/a_192_298#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_75/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_58/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_36/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_75/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_36/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_40/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_24/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_dummy_3v1024x8m81_42/m2_346_89#
+ 018SRAM_cell1_2x_3v1024x8m81_24/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_40/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_39/a_192_298# 018SRAM_cell1_dummy_R_3v1024x8m81_73/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_56/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_3v1024x8m81_42/m2_134_89#
+ 018SRAM_cell1_2x_3v1024x8m81_56/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_50/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_12/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v1024x8m81_85/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_46/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_85/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_46/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_dummy_3v1024x8m81_4/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_52/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_13/m2_346_89# 018SRAM_cell1_2x_3v1024x8m81_54/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_4/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_52/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_13/m2_134_89# 018SRAM_cell1_2x_3v1024x8m81_54/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_101/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_25/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_101/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_58/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_25/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_95/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_17/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_56/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_35/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_95/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_56/a_248_342# 018SRAM_cell1_dummy_3v1024x8m81_62/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_17/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_41/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_3v1024x8m81_23/m2_346_89# 018SRAM_cell1_dummy_R_3v1024x8m81_59/a_192_298#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_111/m3_82_330# 018SRAM_cell1_dummy_3v1024x8m81_23/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_62/m2_134_89# 018SRAM_cell1_2x_3v1024x8m81_57/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_111/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_66/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_39/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_27/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_39/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_54/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_27/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_87/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_66/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_40/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_3v1024x8m81_33/m2_346_89# 018SRAM_cell1_dummy_R_3v1024x8m81_69/a_192_298#
+ 018SRAM_cell1_dummy_3v1024x8m81_33/m2_134_89# 018SRAM_cell1_dummy_R_3v1024x8m81_121/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_121/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_25/018SRAM_cell1_3v1024x8m81_1/a_248_592# 018SRAM_cell1_2x_3v1024x8m81_53/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_76/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_37/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_53/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_76/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_24/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_37/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_43/m2_346_89# 018SRAM_cell1_dummy_R_3v1024x8m81_79/a_192_298#
+ 018SRAM_cell1_2x_3v1024x8m81_24/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_83/w_30_512#
+ 018SRAM_cell1_dummy_3v1024x8m81_43/m2_134_89# 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_39/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_86/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_56/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_47/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_86/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_47/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_22/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_5/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_53/m2_346_89#
+ 018SRAM_cell1_2x_3v1024x8m81_22/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_89/a_192_298#
+ 018SRAM_cell1_dummy_3v1024x8m81_14/m2_346_89# 018SRAM_cell1_2x_3v1024x8m81_38/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_54/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_5/m2_134_89# 018SRAM_cell1_dummy_R_3v1024x8m81_102/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_54/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_38/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_3v1024x8m81_14/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_53/m2_134_89# 018SRAM_cell1_2x_3v1024x8m81_54/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_102/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_35/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_105/a_192_298#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_96/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_57/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_18/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_18/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_96/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_57/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v1024x8m81_18/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_24/m2_346_89# 018SRAM_cell1_dummy_R_3v1024x8m81_99/a_192_298#
+ 018SRAM_cell1_dummy_3v1024x8m81_63/m2_346_89# 018SRAM_cell1_2x_3v1024x8m81_52/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_0/a_192_298# 018SRAM_cell1_dummy_3v1024x8m81_63/m2_134_89#
+ 018SRAM_cell1_2x_3v1024x8m81_52/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_112/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_24/m2_134_89# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_112/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_59/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_115/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_39/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_67/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_31/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_28/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_39/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_67/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_28/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_97/w_30_512# 018SRAM_cell1_dummy_3v1024x8m81_34/m2_346_89#
+ m3_15667_n5552# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_3v1024x8m81_34/m2_134_89# 018SRAM_cell1_dummy_R_3v1024x8m81_122/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_21/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_21/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_122/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_37/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_53/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_125/a_192_298# 018SRAM_cell1_dummy_R_3v1024x8m81_109/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_77/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_38/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_53/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_37/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_38/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_77/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_44/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_dummy_3v1024x8m81_44/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_60/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_93/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_7/w_30_512# 018SRAM_cell1_dummy_3v1024x8m81_44/m2_134_89#
+ 018SRAM_cell1_2x_3v1024x8m81_32/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_2x_3v1024x8m81_51/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_40/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v1024x8m81_48/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_248_592# ypass_gate_3v1024x8m81_0_0/vdd_uq0
+ 018SRAM_cell1_dummy_R_3v1024x8m81_87/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_51/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_87/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_22/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_48/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_105/w_30_512#
+ 018SRAM_cell1_dummy_3v1024x8m81_6/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_54/m2_346_89#
+ 018SRAM_cell1_2x_3v1024x8m81_22/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_3v1024x8m81_15/m2_346_89# 018SRAM_cell1_dummy_R_3v1024x8m81_40/a_192_298#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_38/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_54/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_6/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_15/m2_134_89# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_38/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_103/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_8/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_103/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_97/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_54/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_58/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_20/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_58/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_97/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_64/m2_346_89# 018SRAM_cell1_2x_3v1024x8m81_20/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_25/m2_346_89# 018SRAM_cell1_dummy_R_3v1024x8m81_1/a_192_298#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_36/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_52/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_101/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_36/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_3v1024x8m81_64/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_113/m3_82_330# 018SRAM_cell1_dummy_3v1024x8m81_25/m2_134_89#
+ 018SRAM_cell1_2x_3v1024x8m81_52/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_34/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_15667_n6510#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_113/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_2/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_2/a_248_342# pmos_5p04310591302095_3v1024x8m81_0/S
+ 018SRAM_cell1_dummy_R_3v1024x8m81_68/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_29/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_64/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_29/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_68/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_35/m2_346_89# 018SRAM_cell1_dummy_R_3v1024x8m81_60/a_192_298#
+ 018SRAM_cell1_2x_3v1024x8m81_50/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_39/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_50/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_dummy_3v1024x8m81_35/m2_134_89# 018SRAM_cell1_dummy_R_3v1024x8m81_123/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_21/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_123/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_21/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_39/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_37/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_119/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_39/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_37/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_78/m3_82_330#
+ ypass_gate_3v1024x8m81_0_0/vdd 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_78/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_39/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_45/m2_346_89# 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_31/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_53/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_3v1024x8m81_45/m2_134_89# 018SRAM_cell1_dummy_R_3v1024x8m81_59/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_35/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ m3_15667_n6288# 018SRAM_cell1_2x_3v1024x8m81_51/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_88/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_51/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_35/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_49/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_32/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_88/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_115/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_49/a_248_342# 018SRAM_cell1_dummy_3v1024x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_55/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_16/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_64/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_3v1024x8m81_55/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_7/m2_134_89#
+ 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v1024x8m81_104/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_16/m2_134_89# 018SRAM_cell1_dummy_R_3v1024x8m81_104/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_55/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_38/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v1024x8m81_59/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_98/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_107/a_192_298#
+ 018SRAM_cell1_2x_3v1024x8m81_20/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_98/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_59/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_53/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_20/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_26/m2_346_89# 018SRAM_cell1_2x_3v1024x8m81_36/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_111/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_8/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_36/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v1024x8m81_26/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_114/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_3/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_114/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_52/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_3/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_117/a_192_298#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_69/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_69/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_36/m2_346_89# 018SRAM_cell1_2x_3v1024x8m81_34/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_50/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_61/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_58/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_50/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_34/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_13/018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_124/m3_82_330# 018SRAM_cell1_dummy_3v1024x8m81_36/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_124/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_79/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_127/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_79/a_248_342# m3_15698_n15942# 018SRAM_cell1_dummy_3v1024x8m81_46/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_71/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_37/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_32/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_36/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_69/w_30_512#
+ 018SRAM_cell1_dummy_3v1024x8m81_46/m2_134_89# m2_16574_21# 018SRAM_cell1_2x_3v1024x8m81_43/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_35/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_89/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_35/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_89/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_125/w_30_512#
+ 018SRAM_cell1_dummy_3v1024x8m81_56/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_81/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_51/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_3v1024x8m81_17/m2_346_89# m3_15667_n7247# 018SRAM_cell1_dummy_3v1024x8m81_8/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_56/m2_134_89# 018SRAM_cell1_dummy_R_3v1024x8m81_105/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_17/m2_134_89# 018SRAM_cell1_dummy_R_3v1024x8m81_32/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_65/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_105/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_3/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_3/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_99/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_10/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_99/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_60/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_10/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_91/a_192_298#
+ 018SRAM_cell1_dummy_3v1024x8m81_27/m2_346_89# 018SRAM_cell1_dummy_R_3v1024x8m81_6/a_192_298#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_121/w_30_512# 018SRAM_cell1_dummy_3v1024x8m81_27/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_115/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_4/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_115/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_4/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_36/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_63/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_20/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_61/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_5/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_20/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_63/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_18/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_dummy_3v1024x8m81_37/m2_346_89#
+ 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_62/a_192_298#
+ 018SRAM_cell1_2x_3v1024x8m81_34/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_18/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_34/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_37/m2_134_89# 018SRAM_cell1_dummy_R_3v1024x8m81_125/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_125/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_30/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_30/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_32/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_dummy_3v1024x8m81_47/m2_346_89#
+ 018SRAM_cell1_2x_3v1024x8m81_2/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_2/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_38/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_32/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_33/a_192_298#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_6/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_48/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_47/m2_134_89# 018SRAM_cell1_dummy_R_3v1024x8m81_79/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_48/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_63/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v1024x8m81_40/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_40/a_248_342# pmos_5p04310591302097_3v1024x8m81_0/S
+ 018SRAM_cell1_dummy_3v1024x8m81_18/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_57/m2_346_89#
+ 018SRAM_cell1_2x_3v1024x8m81_35/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_dummy_3v1024x8m81_9/m2_346_89#
+ 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_1/a_248_592# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_57/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_9/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_18/m2_134_89# 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_106/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_53/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_106/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_3/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_75/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_3/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_50/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_109/a_192_298#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_11/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_11/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_50/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v1024x8m81_28/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_53/a_192_298# 018SRAM_cell1_dummy_R_3v1024x8m81_2/a_192_298#
+ m3_15645_n13711# 018SRAM_cell1_2x_3v1024x8m81_48/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_116/m3_82_330# 018SRAM_cell1_dummy_3v1024x8m81_28/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_5/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_1/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_31/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_116/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_31/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_5/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_52/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_1/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_119/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_47/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_63/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_71/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_60/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_21/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_47/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_60/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_63/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_21/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_18/018SRAM_cell1_3v1024x8m81_1/m3_82_330# ypass_gate_3v1024x8m81_0_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ 018SRAM_cell1_dummy_3v1024x8m81_38/m2_346_89# 018SRAM_cell1_dummy_R_3v1024x8m81_63/a_192_298#
+ 018SRAM_cell1_2x_3v1024x8m81_18/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v1024x8m81_38/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_126/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_34/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_126/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_3/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_61/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_70/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_57/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_50/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_61/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_31/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_70/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_31/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_32/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_16/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_2/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_16/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_45/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_73/a_192_298# 018SRAM_cell1_dummy_3v1024x8m81_48/m2_346_89#
+ 018SRAM_cell1_2x_3v1024x8m81_2/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_34/a_192_298#
+ 018SRAM_cell1_2x_3v1024x8m81_32/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_56/w_30_512#
+ 018SRAM_cell1_dummy_3v1024x8m81_48/m2_134_89# 018SRAM_cell1_dummy_R_3v1024x8m81_89/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_48/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_48/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_80/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_41/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_80/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_0/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_41/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_42/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_dummy_3v1024x8m81_19/m2_346_89#
+ 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_0/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_83/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_19/m2_134_89# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_107/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_107/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_85/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_90/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_51/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_12/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_90/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_51/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v1024x8m81_12/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_29/m2_346_89# 018SRAM_cell1_dummy_R_3v1024x8m81_93/a_192_298#
+ 018SRAM_cell1_2x_3v1024x8m81_60/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_54/a_192_298#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_4/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_47/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_60/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_117/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_15/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_29/m2_134_89# 018SRAM_cell1_2x_3v1024x8m81_31/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_117/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_1/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_6/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_31/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_15/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_6/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_1/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_47/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_61/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_81/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_22/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_61/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_22/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_47/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_37/w_30_512# 018SRAM_cell1_dummy_3v1024x8m81_39/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_127/m3_82_330# 018SRAM_cell1_dummy_3v1024x8m81_39/m2_134_89#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_31/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_127/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_45/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_61/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_71/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_32/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_61/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_45/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_71/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_16/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_32/a_248_342# 018SRAM_cell1_dummy_3v1024x8m81_49/m2_346_89#
+ 018SRAM_cell1_2x_3v1024x8m81_16/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_35/a_192_298#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_33/w_30_512# 018SRAM_cell1_dummy_3v1024x8m81_49/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_99/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_31/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_0/a_248_592# m3_15667_n6043#
+ 018SRAM_cell1_2x_3v1024x8m81_61/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_37/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_81/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_42/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_42/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_14/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_81/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_0/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_3v1024x8m81_0/m2_346_89#
+ 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_14/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_59/m2_346_89# 018SRAM_cell1_2x_3v1024x8m81_0/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_3v1024x8m81_59/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_0/m2_134_89# 018SRAM_cell1_dummy_R_3v1024x8m81_108/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_62/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_95/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_108/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_3/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_91/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_52/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_13/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_91/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_52/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v1024x8m81_13/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_55/a_192_298#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_7/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_44/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_60/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_44/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_60/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_118/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_107/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_15/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_7/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_118/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_7/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_15/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_62/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_23/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_62/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_91/w_30_512# 018SRAM_cell1_dummy_R_3v1024x8m81_2/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_1/a_248_592# 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_23/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_65/a_192_298#
+ 018SRAM_cell1_2x_3v1024x8m81_51/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_47/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_13/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_13/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_103/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_45/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_72/m3_82_330#
+ ypass_gate_3v1024x8m81_0_0/pcb 018SRAM_cell1_dummy_R_3v1024x8m81_33/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_45/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_72/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_33/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_75/a_192_298#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_36/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_61/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_0/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_56/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_18/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_2x_3v1024x8m81_11/018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_43/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_43/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_43/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_82/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_82/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_14/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_59/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_43/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_1/m2_346_89# 018SRAM_cell1_2x_3v1024x8m81_59/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_14/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v1024x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_85/a_192_298# m3_15667_n7002# 018SRAM_cell1_dummy_3v1024x8m81_1/m2_134_89#
+ m2_16574_77581# 018SRAM_cell1_dummy_R_3v1024x8m81_109/m3_82_330# 018SRAM_cell1_dummy_3v1024x8m81_10/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_109/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_40/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_2x_3v1024x8m81_41/018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_101/a_192_298# 018SRAM_cell1_dummy_R_3v1024x8m81_92/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v1024x8m81_53/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_14/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_12/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_53/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_92/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_12/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_14/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_20/m2_346_89# 018SRAM_cell1_dummy_R_3v1024x8m81_95/a_192_298#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_5/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_44/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_56/a_192_298# 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ a_n547_178# 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_44/018SRAM_cell1_3v1024x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_117/w_30_512#
+ VSUBS 018SRAM_cell1_dummy_3v1024x8m81_20/m2_134_89# 018SRAM_cell1_dummy_R_3v1024x8m81_119/m3_82_330#
+ m3_n631_83# 018SRAM_cell1_dummy_R_3v1024x8m81_8/m3_82_330# 018SRAM_cell1_dummy_R_3v1024x8m81_119/a_248_342#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_8/a_248_342# 018SRAM_cell1_dummy_R_3v1024x8m81_63/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_111/a_192_298# 018SRAM_cell1_dummy_R_3v1024x8m81_24/m3_82_330#
+ m3_15667_n6752# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_0/w_30_512#
X018SRAM_cell1_3v1024x8m81_1 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ m3_n631_83# 018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# VSUBS x018SRAM_cell1_3v1024x8m81
Xpmos_5p04310591302095_3v1024x8m81_0 pmos_5p04310591302095_3v1024x8m81_0/D ypass_gate_3v1024x8m81_0_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_0_0/pmos_5p0431059130201_3v1024x8m81_0/D pmos_5p04310591302095_3v1024x8m81_0/S
+ pmos_5p04310591302095_3v1024x8m81_0/S pmos_5p04310591302095_3v1024x8m81_0/S pmos_5p04310591302095_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_90 018SRAM_cell1_dummy_R_3v1024x8m81_90/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_90/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_91/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_91/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_60 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_60/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_60/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_80 018SRAM_cell1_dummy_R_3v1024x8m81_80/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_80/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_81/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_81/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_91 018SRAM_cell1_dummy_R_3v1024x8m81_91/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_91/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_91/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_91/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_120 018SRAM_cell1_dummy_R_3v1024x8m81_120/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_120/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_121/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_121/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_61 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_61/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_61/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_50 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_50/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_50/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_92 018SRAM_cell1_dummy_R_3v1024x8m81_92/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_92/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_93/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_93/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_70 018SRAM_cell1_dummy_R_3v1024x8m81_70/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_70/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_71/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_71/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_81 018SRAM_cell1_dummy_R_3v1024x8m81_81/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_81/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_81/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_81/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_121 018SRAM_cell1_dummy_R_3v1024x8m81_121/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_121/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_121/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_121/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_110 018SRAM_cell1_dummy_R_3v1024x8m81_110/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_110/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_111/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_111/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_62 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_62/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_62/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_51 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_51/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_51/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_40 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_40/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_40/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_93 018SRAM_cell1_dummy_R_3v1024x8m81_93/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_93/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_93/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_93/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_60 018SRAM_cell1_dummy_R_3v1024x8m81_60/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_60/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_60/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_60/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_71 018SRAM_cell1_dummy_R_3v1024x8m81_71/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_71/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_71/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_71/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_82 018SRAM_cell1_dummy_R_3v1024x8m81_82/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_82/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_83/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_83/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_122 018SRAM_cell1_dummy_R_3v1024x8m81_122/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_122/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_123/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_123/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_111 018SRAM_cell1_dummy_R_3v1024x8m81_111/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_111/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_111/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_111/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_100 018SRAM_cell1_dummy_R_3v1024x8m81_100/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_100/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_101/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_101/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_63 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_63/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_63/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_52 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_52/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_52/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_41 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_41/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_41/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_30 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_30/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_30/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_94 018SRAM_cell1_dummy_R_3v1024x8m81_94/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_94/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_95/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_95/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_50 018SRAM_cell1_dummy_R_3v1024x8m81_50/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_50/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_60/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_60/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_61 018SRAM_cell1_dummy_R_3v1024x8m81_61/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_61/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_61/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_61/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_72 018SRAM_cell1_dummy_R_3v1024x8m81_72/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_72/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_73/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_73/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_83 018SRAM_cell1_dummy_R_3v1024x8m81_83/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_83/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_83/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_83/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_123 018SRAM_cell1_dummy_R_3v1024x8m81_123/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_123/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_123/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_123/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_112 018SRAM_cell1_dummy_R_3v1024x8m81_112/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_112/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_113/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_113/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_101 018SRAM_cell1_dummy_R_3v1024x8m81_101/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_101/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_101/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_101/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_64 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_64/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_64/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_53 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_53/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_53/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_42 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_42/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_42/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_20 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_20/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_20/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_31 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_31/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_31/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_95 018SRAM_cell1_dummy_R_3v1024x8m81_95/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_95/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_95/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_95/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_40 018SRAM_cell1_dummy_R_3v1024x8m81_40/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_40/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_40/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_40/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_62 018SRAM_cell1_dummy_R_3v1024x8m81_62/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_62/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_62/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_62/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_51 018SRAM_cell1_dummy_R_3v1024x8m81_51/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_51/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_58/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_58/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_73 018SRAM_cell1_dummy_R_3v1024x8m81_73/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_73/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_73/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_73/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_84 018SRAM_cell1_dummy_R_3v1024x8m81_84/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_84/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_85/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_85/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_124 018SRAM_cell1_dummy_R_3v1024x8m81_124/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_124/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_125/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_125/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_113 018SRAM_cell1_dummy_R_3v1024x8m81_113/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_113/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_113/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_113/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_102 018SRAM_cell1_dummy_R_3v1024x8m81_102/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_102/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_103/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_103/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_54 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_54/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_54/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_43 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_43/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_43/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_32 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_32/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_32/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_10 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_10/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_21 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_21/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_21/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
Xpmos_5p04310591302097_3v1024x8m81_0 pmos_5p04310591302097_3v1024x8m81_0/D pmos_5p04310591302095_3v1024x8m81_0/D
+ pmos_5p04310591302095_3v1024x8m81_0/D w_15880_n13729# pmos_5p04310591302097_3v1024x8m81_0/S
+ pmos_5p04310591302097_3v1024x8m81_0/S pmos_5p04310591302097_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_96 018SRAM_cell1_dummy_R_3v1024x8m81_96/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_96/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_97/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_97/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_30 018SRAM_cell1_dummy_R_3v1024x8m81_30/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_30/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_39/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_39/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_41 018SRAM_cell1_dummy_R_3v1024x8m81_41/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_41/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_64/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_64/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_63 018SRAM_cell1_dummy_R_3v1024x8m81_63/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_63/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_63/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_63/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_52 018SRAM_cell1_dummy_R_3v1024x8m81_52/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_52/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_59/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_59/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_74 018SRAM_cell1_dummy_R_3v1024x8m81_74/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_74/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_75/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_75/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_85 018SRAM_cell1_dummy_R_3v1024x8m81_85/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_85/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_85/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_85/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_125 018SRAM_cell1_dummy_R_3v1024x8m81_125/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_125/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_125/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_125/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_114 018SRAM_cell1_dummy_R_3v1024x8m81_114/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_114/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_115/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_115/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_103 018SRAM_cell1_dummy_R_3v1024x8m81_103/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_103/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_103/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_103/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_55 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_55/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_55/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_44 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_44/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_44/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_33 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_33/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_33/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_11 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_11/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_22 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_22/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_22/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_0/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_0/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_0/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_0/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_97 018SRAM_cell1_dummy_R_3v1024x8m81_97/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_97/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_97/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_97/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_31 018SRAM_cell1_dummy_R_3v1024x8m81_31/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_31/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_31/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_31/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_20 018SRAM_cell1_dummy_R_3v1024x8m81_20/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_20/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_31/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_31/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_64 018SRAM_cell1_dummy_R_3v1024x8m81_64/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_64/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_64/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_64/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_53 018SRAM_cell1_dummy_R_3v1024x8m81_53/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_53/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_53/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_53/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_42 018SRAM_cell1_dummy_R_3v1024x8m81_42/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_42/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_53/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_53/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_75 018SRAM_cell1_dummy_R_3v1024x8m81_75/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_75/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_75/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_75/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_86 018SRAM_cell1_dummy_R_3v1024x8m81_86/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_86/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_87/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_87/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_126 018SRAM_cell1_dummy_R_3v1024x8m81_126/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_126/a_248_342# m2_16574_77581# 018SRAM_cell1_dummy_R_3v1024x8m81_127/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_127/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_115 018SRAM_cell1_dummy_R_3v1024x8m81_115/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_115/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_115/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_115/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_104 018SRAM_cell1_dummy_R_3v1024x8m81_104/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_104/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_105/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_105/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_56 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_56/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_56/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_45 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_45/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_45/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_34 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_34/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_34/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_1/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_1/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_1/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_1/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_12 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_12/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_23 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_23/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_23/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_98 018SRAM_cell1_dummy_R_3v1024x8m81_98/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_98/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_99/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_99/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_10 018SRAM_cell1_dummy_R_3v1024x8m81_10/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_10/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_0/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_0/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_65 018SRAM_cell1_dummy_R_3v1024x8m81_65/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_65/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_65/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_65/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_21 018SRAM_cell1_dummy_R_3v1024x8m81_21/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_21/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_35/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_35/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_32 018SRAM_cell1_dummy_R_3v1024x8m81_32/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_32/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_32/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_32/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_54 018SRAM_cell1_dummy_R_3v1024x8m81_54/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_54/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_54/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_54/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_43 018SRAM_cell1_dummy_R_3v1024x8m81_43/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_43/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_57/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_57/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_76 018SRAM_cell1_dummy_R_3v1024x8m81_76/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_76/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_77/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_77/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_87 018SRAM_cell1_dummy_R_3v1024x8m81_87/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_87/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_87/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_87/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_127 018SRAM_cell1_dummy_R_3v1024x8m81_127/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_127/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_127/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_127/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_116 018SRAM_cell1_dummy_R_3v1024x8m81_116/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_116/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_117/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_117/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_105 018SRAM_cell1_dummy_R_3v1024x8m81_105/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_105/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_105/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_105/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_57 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_57/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_57/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_46 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_46/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_46/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_35 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_35/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_35/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_2/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_2/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_2/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_2/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_13 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_13/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_24 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_24/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_24/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_99 018SRAM_cell1_dummy_R_3v1024x8m81_99/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_99/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_99/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_99/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_11 018SRAM_cell1_dummy_R_3v1024x8m81_11/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_11/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_1/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_1/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_33 018SRAM_cell1_dummy_R_3v1024x8m81_33/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_33/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_33/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_33/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_22 018SRAM_cell1_dummy_R_3v1024x8m81_22/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_22/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_37/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_37/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_55 018SRAM_cell1_dummy_R_3v1024x8m81_55/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_55/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_55/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_55/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_44 018SRAM_cell1_dummy_R_3v1024x8m81_44/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_44/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_55/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_55/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_66 018SRAM_cell1_dummy_R_3v1024x8m81_66/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_66/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_67/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_67/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_77 018SRAM_cell1_dummy_R_3v1024x8m81_77/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_77/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_77/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_77/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_88 018SRAM_cell1_dummy_R_3v1024x8m81_88/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_88/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_89/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_89/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_128 m2_16574_77581# VSUBS m2_16574_77581# 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_117 018SRAM_cell1_dummy_R_3v1024x8m81_117/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_117/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_117/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_117/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_106 018SRAM_cell1_dummy_R_3v1024x8m81_106/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_106/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_107/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_107/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_47 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_47/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_47/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_36 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_36/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_36/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_14 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_14/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_25 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_25/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_25/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_3/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_3/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_3/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_3/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_3/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_3/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_12 018SRAM_cell1_dummy_R_3v1024x8m81_12/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_12/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_8/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_8/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_34 018SRAM_cell1_dummy_R_3v1024x8m81_34/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_34/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_34/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_34/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_23 018SRAM_cell1_dummy_R_3v1024x8m81_23/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_23/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_36/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_36/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_45 018SRAM_cell1_dummy_R_3v1024x8m81_45/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_45/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_62/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_62/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_56 018SRAM_cell1_dummy_R_3v1024x8m81_56/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_56/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_56/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_56/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_67 018SRAM_cell1_dummy_R_3v1024x8m81_67/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_67/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_67/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_67/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_78 018SRAM_cell1_dummy_R_3v1024x8m81_78/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_78/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_79/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_79/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_89 018SRAM_cell1_dummy_R_3v1024x8m81_89/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_89/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_89/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_89/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_129 018SRAM_cell1_dummy_R_3v1024x8m81_129/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_129/a_248_342# m2_16574_77581# 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_118 018SRAM_cell1_dummy_R_3v1024x8m81_118/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_118/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_119/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_119/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_107 018SRAM_cell1_dummy_R_3v1024x8m81_107/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_107/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_107/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_107/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_59 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_59/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_59/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_48 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_48/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_48/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_37 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_37/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_37/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_4 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_4/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_15 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_15/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_26 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_26/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_26/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_13 018SRAM_cell1_dummy_R_3v1024x8m81_13/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_13/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_6/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_6/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_35 018SRAM_cell1_dummy_R_3v1024x8m81_35/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_35/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_35/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_35/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_24 018SRAM_cell1_dummy_R_3v1024x8m81_24/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_24/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_32/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_32/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_46 018SRAM_cell1_dummy_R_3v1024x8m81_46/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_46/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_54/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_54/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_57 018SRAM_cell1_dummy_R_3v1024x8m81_57/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_57/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_57/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_57/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_68 018SRAM_cell1_dummy_R_3v1024x8m81_68/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_68/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_69/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_69/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_79 018SRAM_cell1_dummy_R_3v1024x8m81_79/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_79/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_79/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_79/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_119 018SRAM_cell1_dummy_R_3v1024x8m81_119/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_119/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_119/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_119/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_108 018SRAM_cell1_dummy_R_3v1024x8m81_108/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_108/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_109/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_109/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_49 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_49/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_49/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_38 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_38/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_38/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_16 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_16/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_16/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_27 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_27/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_27/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_5 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_5/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
Xnmos_5p04310591302096_3v1024x8m81_0 pmos_5p04310591302097_3v1024x8m81_0/D pmos_5p04310591302095_3v1024x8m81_0/D
+ pmos_5p04310591302095_3v1024x8m81_0/D VSUBS VSUBS VSUBS nmos_5p04310591302096_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_14 018SRAM_cell1_dummy_R_3v1024x8m81_14/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_14/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_2/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_2/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_25 018SRAM_cell1_dummy_R_3v1024x8m81_25/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_25/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_33/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_33/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_36 018SRAM_cell1_dummy_R_3v1024x8m81_36/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_36/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_36/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_36/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_58 018SRAM_cell1_dummy_R_3v1024x8m81_58/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_58/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_58/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_58/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_47 018SRAM_cell1_dummy_R_3v1024x8m81_47/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_47/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_56/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_56/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_69 018SRAM_cell1_dummy_R_3v1024x8m81_69/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_69/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_69/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_69/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_60 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_61/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_60/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_61/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_60/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_60/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_60/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_60/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_60/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_0 018SRAM_cell1_dummy_R_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_0/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_0/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_0/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_109 018SRAM_cell1_dummy_R_3v1024x8m81_109/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_109/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_109/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_109/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_39 m2_16574_77581# VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# m2_16574_77581# 018SRAM_cell1_dummy_3v1024x8m81_39/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_39/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_6 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_6/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_17 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_17/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_17/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_28 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_28/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_28/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_15 018SRAM_cell1_dummy_R_3v1024x8m81_15/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_15/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_4/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_4/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_26 018SRAM_cell1_dummy_R_3v1024x8m81_26/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_26/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_65/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_65/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_37 018SRAM_cell1_dummy_R_3v1024x8m81_37/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_37/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_37/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_37/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_48 018SRAM_cell1_dummy_R_3v1024x8m81_48/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_48/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_61/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_61/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_59 018SRAM_cell1_dummy_R_3v1024x8m81_59/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_59/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_59/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_59/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_61 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_61/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_61/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_61/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_61/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_61/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_61/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_50 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_51/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_50/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_51/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_50/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_50/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_50/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_50/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_50/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_1 018SRAM_cell1_dummy_R_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_1/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_1/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_1/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
Xypass_gate_3v1024x8m81_0_0 ypass_gate_3v1024x8m81_0_0/vss ypass_gate_3v1024x8m81_0_0/bb
+ ypass_gate_3v1024x8m81_0_0/db ypass_gate_3v1024x8m81_0_0/ypass ypass_gate_3v1024x8m81_0_0/d
+ ypass_gate_3v1024x8m81_0_0/pcb ypass_gate_3v1024x8m81_0_0/vdd_uq0 m3_15667_n7247#
+ ypass_gate_3v1024x8m81_0_0/bb m3_15667_n6510# ypass_gate_3v1024x8m81_0_0/vdd_uq0
+ m3_15667_n6288# ypass_gate_3v1024x8m81_0_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ m3_15667_n5552# ypass_gate_3v1024x8m81_0_0/vdd_uq0 VSUBS m3_15667_n5798# ypass_gate_3v1024x8m81_0_0/b
+ m3_15667_n6043# m3_15667_n7002# ypass_gate_3v1024x8m81_0_0/vdd m3_15667_n6752# ypass_gate_3v1024x8m81_0
X018SRAM_cell1_2x_3v1024x8m81_7 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_7/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_18 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_18/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_18/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_29 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_29/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_29/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_16 018SRAM_cell1_dummy_R_3v1024x8m81_16/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_16/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_7/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_7/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_38 018SRAM_cell1_dummy_R_3v1024x8m81_38/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_38/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_38/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_38/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_27 018SRAM_cell1_dummy_R_3v1024x8m81_27/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_27/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_38/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_38/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_49 018SRAM_cell1_dummy_R_3v1024x8m81_49/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_49/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_63/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_63/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_62 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_63/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_63/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_62/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_51 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_52/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_51/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_52/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_51/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_51/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_51/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_51/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_51/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_40 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_41/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_40/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_41/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_40/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_40/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_40/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_40/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_40/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_2 018SRAM_cell1_dummy_R_3v1024x8m81_2/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_2/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_2/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_2/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_8 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_8/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_19 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_19/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_19/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_17 018SRAM_cell1_dummy_R_3v1024x8m81_17/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_17/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_5/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_5/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_39 018SRAM_cell1_dummy_R_3v1024x8m81_39/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_39/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_39/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_39/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_28 018SRAM_cell1_dummy_R_3v1024x8m81_28/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_28/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_40/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_40/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_63 m3_n631_83# 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v1024x8m81_63/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v1024x8m81_63/018SRAM_cell1_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_63/018SRAM_cell1_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v1024x8m81_63/018SRAM_cell1_3v1024x8m81_0/a_248_592# 018SRAM_cell1_2x_3v1024x8m81_63/018SRAM_cell1_3v1024x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_63/018SRAM_cell1_3v1024x8m81_1/a_248_342# VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_52 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_53/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_52/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_53/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_52/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_52/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_52/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_52/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_52/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_30 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_41 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_42/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_41/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_42/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_41/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_41/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_41/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_41/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_41/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_3 018SRAM_cell1_dummy_R_3v1024x8m81_3/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_3/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_3/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_3/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_9 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_0 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_0/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_18 018SRAM_cell1_dummy_R_3v1024x8m81_18/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_18/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_3/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_3/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_29 018SRAM_cell1_dummy_R_3v1024x8m81_29/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_29/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_34/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_34/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_53 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_54/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_53/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_54/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_53/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_53/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_53/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_53/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_53/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_31 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_31/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_3/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_31/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_31/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_31/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_3/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_31/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_31/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_20 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_25/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_20/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_20/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_25/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_20/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_20/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_42 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_43/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_42/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_43/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_42/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_42/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_42/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_42/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_42/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_4 018SRAM_cell1_dummy_R_3v1024x8m81_4/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_4/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_4/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_4/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_1 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_1/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_19 a_n547_178# VSUBS m2_16574_21# 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_54 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_54/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_54/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_54/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_54/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_54/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_54/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_10 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_12/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_11/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_12/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_10/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_10/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_11/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_10/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_10/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_21 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_21/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_21/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_21/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_21/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_32 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_32/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_32/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_32/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_32/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_32/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_32/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_43 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_44/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_43/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_44/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_43/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_43/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_43/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_43/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_43/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_5 018SRAM_cell1_dummy_R_3v1024x8m81_5/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_5/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_5/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_5/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_2 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_2/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_55 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_56/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_56/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_55/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_11 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_11/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_13/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_11/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_11/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_11/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_13/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_11/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_11/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_22 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_22/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_22/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_22/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_22/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_33 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_34/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_34/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_33/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_44 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_45/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_44/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_45/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_44/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_44/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_44/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_44/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_44/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_6 018SRAM_cell1_dummy_R_3v1024x8m81_6/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_6/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_6/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_6/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_3 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_3/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_56 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_57/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_56/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_57/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_56/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_56/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_56/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_56/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_56/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_45 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_45/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_45/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_45/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_45/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_45/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_45/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_12 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_12/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_12/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_12/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_12/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_12/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_12/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_23 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_32/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_32/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_23/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_34 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_35/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_34/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_35/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_34/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_34/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_34/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_34/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_34/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_7 018SRAM_cell1_dummy_R_3v1024x8m81_7/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_7/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_7/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_7/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_4 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_4/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_57 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_58/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_57/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_58/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_57/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_57/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_57/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_57/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_57/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_46 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_47/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_47/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_46/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_13 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_13/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_13/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_13/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_13/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_13/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_13/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_24 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_24/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_24/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_24/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_24/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_35 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_36/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_35/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_36/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_35/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_35/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_35/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_35/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_35/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_8 018SRAM_cell1_dummy_R_3v1024x8m81_8/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_8/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v1024x8m81_8/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_dummy_R_3v1024x8m81_8/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_5 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_5/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_14 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_31/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_14/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_14/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_31/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_14/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_14/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_58 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_59/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_58/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_59/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_58/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_58/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_58/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_58/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_58/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_47 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_48/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_47/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_48/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_47/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_47/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_47/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_47/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_47/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_25 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_25/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_25/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_25/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_25/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_30/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_25/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_25/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_36 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_37/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_36/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_37/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_36/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_36/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_36/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_36/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_36/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_R_3v1024x8m81_9 018SRAM_cell1_dummy_R_3v1024x8m81_9/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v1024x8m81_9/a_248_342# m2_16574_21# 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ ypass_gate_3v1024x8m81_0_0/bb ypass_gate_3v1024x8m81_0_0/b 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ VSUBS x018SRAM_cell1_dummy_R_3v1024x8m81
Xnmos_5p04310591302098_3v1024x8m81_0 pmos_5p04310591302095_3v1024x8m81_0/D ypass_gate_3v1024x8m81_0_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ ypass_gate_3v1024x8m81_0_0/pmos_5p0431059130201_3v1024x8m81_0/D VSUBS VSUBS VSUBS
+ nmos_5p04310591302098_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_6 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_6/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_59 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_60/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_59/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_60/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_59/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_59/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_59/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_59/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_59/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_48 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_48/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_48/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_48/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_48/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_48/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_48/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_15 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_18/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_18/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_15/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_15/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_15/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_15/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_26 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_26/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_37 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_38/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_37/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_38/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_37/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_37/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_37/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_37/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_37/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_7 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_7/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_49 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_50/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_50/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_49/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_16 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_1/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_16/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_16/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_16/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_16/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_27 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_27/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_38 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_39/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_38/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_39/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_38/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_38/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_38/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_38/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_38/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_8 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_8/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_17 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_17/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_28 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_28/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_39 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_40/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_39/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_40/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_39/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_39/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_39/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_39/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_39/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_9 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_3v1024x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v1024x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_9/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_18 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_18/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_9/018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_18/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_18/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_18/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_18/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_18/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_29 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_29/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_19 m3_n631_83# 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_0/w_30_512# m3_n631_83#
+ 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_0/a_248_342# 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v1024x8m81_19/018SRAM_cell1_3v1024x8m81_1/a_248_342#
+ VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_3v1024x8m81_0 a_n547_178# VSUBS 018SRAM_cell1_3v1024x8m81_0/w_30_512#
+ a_n547_178# 018SRAM_cell1_3v1024x8m81_0/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# VSUBS x018SRAM_cell1_3v1024x8m81
.ends

.subckt saout_R_m2_3v1024x8m81 ypass[1] ypass[4] ypass[5] GWEN datain b[0] bb[7] q
+ vss_uq6 vdd_uq0 vdd_uq1 vdd_uq2 vdd_uq4 vdd_uq6 b[1] b[5] bb[6] bb[2] b[7] bb[5]
+ GWE ypass[7] bb[3] WEN bb[0] b[3] sa_3v1024x8m81_0/pcb men_uq0 vdd sacntl_2_3v1024x8m81_0/vdd_uq0
+ b[2] vdd_uq5 vdd_uq3 b[6] bb[4] ypass[3] ypass[2] ypass[6] ypass[0] b[4] mux821_3v1024x8m81_0/ypass_gate_3v1024x8m81_7/vdd_uq0
+ vss bb[1] vdd_uq7
Xdin_3v1024x8m81_0 vss datain men_uq0 sa_3v1024x8m81_0/db sa_3v1024x8m81_0/d sa_3v1024x8m81_0/wep
+ vdd_uq3 vdd_uq5 sa_3v1024x8m81_0/pcb vss din_3v1024x8m81
Xsacntl_2_3v1024x8m81_0 sa_3v1024x8m81_0/pcb sa_3v1024x8m81_0/se sacntl_2_3v1024x8m81_0/pmos_5p04310591302027_3v1024x8m81_1/S_uq0
+ men_uq0 sacntl_2_3v1024x8m81_0/pmos_5p04310591302027_3v1024x8m81_2/S_uq0 vdd_uq0
+ sacntl_2_3v1024x8m81_0/vdd_uq0 vss sacntl_2_3v1024x8m81
Xsa_3v1024x8m81_0 sa_3v1024x8m81_0/qp sa_3v1024x8m81_0/qn sa_3v1024x8m81_0/wep sa_3v1024x8m81_0/se
+ sa_3v1024x8m81_0/pcb sa_3v1024x8m81_0/db vdd_uq5 vdd_uq3 sa_3v1024x8m81_0/d vss
+ sa_3v1024x8m81
Xmux821_3v1024x8m81_0 b[1] bb[1] bb[2] sa_3v1024x8m81_0/db sa_3v1024x8m81_0/d sa_3v1024x8m81_0/db
+ ypass[7] b[6] ypass[6] ypass[4] bb[7] bb[3] ypass[2] sa_3v1024x8m81_0/d b[2] bb[4]
+ ypass[5] ypass[3] b[3] ypass[1] sa_3v1024x8m81_0/d ypass[0] b[0] sa_3v1024x8m81_0/d
+ bb[0] sa_3v1024x8m81_0/d bb[5] bb[6] sa_3v1024x8m81_0/db sa_3v1024x8m81_0/db sa_3v1024x8m81_0/d
+ ypass[3] ypass[7] ypass[2] ypass[0] b[4] mux821_3v1024x8m81_0/ypass_gate_3v1024x8m81_7/vdd_uq0
+ ypass[5] ypass[1] ypass[4] sa_3v1024x8m81_0/d b[7] b[5] vdd_uq7 vss ypass[6] sa_3v1024x8m81_0/d
+ sa_3v1024x8m81_0/pcb mux821_3v1024x8m81
Xwen_wm1_3v1024x8m81_0 GWEN men_uq0 sa_3v1024x8m81_0/wep vdd WEN vss vdd_uq1 wen_wm1_3v1024x8m81
Xoutbuf_oe_3v1024x8m81_0 sa_3v1024x8m81_0/qp sa_3v1024x8m81_0/qn sa_3v1024x8m81_0/se
+ q GWE vss vdd_uq3 outbuf_oe_3v1024x8m81
.ends

.subckt rcol4_1024_3v1024x8m81 WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[48] WL[50]
+ WL[52] WL[54] WL[56] WL[61] WL[51] WL[29] WL[25] WL[24] WL[20] WL[27] WL[30] WL[18]
+ WL[41] WL[15] WL[38] WL[45] WL[43] WL[40] WL[39] WL[31] WL[14] WL[16] WL[17] WL[26]
+ WL[19] WL[58] WL[60] WL[62] WL[53] WL[47] WL[55] WL[12] WL[8] WL[5] WL[10] WL[13]
+ WL[6] tblhl GWE WL[11] din[7] q[5] q[6] q[7] din[5] din[6] q[4] pcb[6] pcb[7] WEN[4]
+ WEN[7] pcb[5] WEN[5] WEN[6] d[4] rarray4_1024_3v1024x8m81_0/m3_n1397_25249# rarray4_1024_3v1024x8m81_0/m3_n1397_42217#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_24535# rarray4_1024_3v1024x8m81_0/m3_n1397_60397#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_41503# rarray4_1024_3v1024x8m81_0/m3_n1397_8779#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_68881# rdummy_3v512x4_3v1024x8m81_0/ypass_gate_3v1024x8m81_0_0/pcb
+ rarray4_1024_3v1024x8m81_0/m3_n1397_57259# rarray4_1024_3v1024x8m81_0/m3_n1397_8281#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_74227# rarray4_1024_3v1024x8m81_0/m3_n1397_48277#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_65245# rarray4_1024_3v1024x8m81_0/m3_n1397_47563#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_64531# rarray4_1024_3v1024x8m81_0/m3_n1397_73729#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_20899# rarray4_1024_3v1024x8m81_0/m3_n1397_10705#
+ WL[0] rarray4_1024_3v1024x8m81_0/m3_n1397_43429# rarray4_1024_3v1024x8m81_0/m3_n1397_70093#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_42715# rarray4_1024_3v1024x8m81_0/m3_n1397_60895#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_50701# rarray4_1024_3v1024x8m81_0/m3_n1397_9493#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_75439# rarray4_1024_3v1024x8m81_0/m3_n1397_13129#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_49489# rarray4_1024_3v1024x8m81_0/m3_n1397_66457#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_48775# rarray4_1024_3v1024x8m81_0/m3_n1397_65743#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_5143# rarray4_1024_3v1024x8m81_0/m3_n1397_39793#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_11917# rarray4_1024_3v1024x8m81_0/m3_n1397_56761#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_45139# rarray4_1024_3v1024x8m81_0/m3_n1397_62107#
+ WL[7] WL[57] rarray4_1024_3v1024x8m81_0/m3_n1397_53125# rarray4_1024_3v1024x8m81_0/m3_n1397_3931#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_35443# rarray4_1024_3v1024x8m81_0/m3_n1397_61609#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_52411# WL[42] rdummy_3v512x4_3v1024x8m81_0/m2_16574_21#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_43927# WL[1] rarray4_1024_3v1024x8m81_0/m3_n1397_70591#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_26461# WL[28] rarray4_1024_3v1024x8m81_0/m3_n1397_51913#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_68167# rarray4_1024_3v1024x8m81_0/m3_n1397_59185#
+ pcb[4] WL[49] rarray4_1024_3v1024x8m81_0/m3_n1397_22111# rarray4_1024_3v1024x8m81_0/m3_n1397_76153#
+ WL[21] rarray4_1024_3v1024x8m81_0/m3_n1397_58471# rarray4_1024_3v1024x8m81_0/m3_n1397_67669#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_40291# rarray4_1024_3v1024x8m81_0/m3_n1397_49987#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_66955# rarray4_1024_3v1024x8m81_0/m3_n1397_6355#
+ rdummy_3v512x4_3v1024x8m81_0/m2_16574_77581# rarray4_1024_3v1024x8m81_0/m3_n1397_57973#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_74941# rarray4_1024_3v1024x8m81_0/m3_n1397_63319#
+ WL[9] WL[59] WL[44] rarray4_1024_3v1024x8m81_0/m3_n1397_54337# rarray4_1024_3v1024x8m81_0/m3_n1397_19687#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_71305# rarray4_1024_3v1024x8m81_0/m3_n1397_36655#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_53623# saout_m2_3v1024x8m81_3/ypass[0] rarray4_1024_3v1024x8m81_0/m3_n1397_27673#
+ saout_R_m2_3v1024x8m81_3/vdd rarray4_1024_3v1024x8m81_0/m3_n1397_44641# WL[2] saout_m2_3v1024x8m81_3/ypass[1]
+ saout_m2_3v1024x8m81_3/VDD_uq0 rarray4_1024_3v1024x8m81_0/m3_n1397_69379# rarray4_1024_3v1024x8m81_0/m3_n1397_51199#
+ saout_m2_3v1024x8m81_3/ypass[2] rarray4_1024_3v1024x8m81_0/m3_n1397_24037# saout_m2_3v1024x8m81_3/vdd_uq2
+ rarray4_1024_3v1024x8m81_0/m3_n1397_41005# rarray4_1024_3v1024x8m81_0/m3_n1397_23323#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_77365# saout_m2_3v1024x8m81_3/ypass[3] WL[23]
+ rarray4_1024_3v1024x8m81_0/m3_n1397_59683# rarray4_1024_3v1024x8m81_0/m3_n1397_76651#
+ WL[22] saout_m2_3v1024x8m81_3/ypass[4] saout_m2_3v1024x8m81_3/men rarray4_1024_3v1024x8m81_0/m3_n1397_7567#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_39079# saout_m2_3v1024x8m81_3/ypass[5] rarray4_1024_3v1024x8m81_0/m3_n1397_56047#
+ saout_m2_3v1024x8m81_3/vdd rarray4_1024_3v1024x8m81_0/m3_n1397_73015# saout_m2_3v1024x8m81_3/vdd_uq0
+ saout_m2_3v1024x8m81_3/ypass[6] rarray4_1024_3v1024x8m81_0/m3_n1397_47065# rarray4_1024_3v1024x8m81_0/m3_n1397_64033#
+ WL[46] rarray4_1024_3v1024x8m81_0/m3_n1397_55549# rarray4_1024_3v1024x8m81_0/m3_n1397_46351#
+ saout_m2_3v1024x8m81_3/ypass[7] rarray4_1024_3v1024x8m81_0/m3_n1397_72517# rarray4_1024_3v1024x8m81_0/m3_n1397_37867#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_54835# saout_m2_3v1024x8m81_3/vdd_uq1 saout_m2_3v1024x8m81_3/GWEN
+ rarray4_1024_3v1024x8m81_0/m3_n1397_71803# rarray4_1024_3v1024x8m81_0/m3_n1397_28885#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_45853# WL[4] saout_m2_3v1024x8m81_3/VDD rarray4_1024_3v1024x8m81_0/m3_n1397_62821#
+ saout_m2_3v1024x8m81_3/vdd_uq3 WL[3] VSS
Xsaout_m2_3v1024x8m81_2 saout_m2_3v1024x8m81_3/ypass[1] saout_m2_3v1024x8m81_3/ypass[2]
+ saout_m2_3v1024x8m81_3/ypass[4] saout_m2_3v1024x8m81_3/ypass[0] saout_m2_3v1024x8m81_3/GWEN
+ din[6] q[6] saout_m2_3v1024x8m81_2/pcb saout_m2_3v1024x8m81_2/bb[0] saout_m2_3v1024x8m81_2/b[0]
+ saout_m2_3v1024x8m81_2/bb[1] saout_m2_3v1024x8m81_2/b[2] saout_m2_3v1024x8m81_2/b[5]
+ saout_m2_3v1024x8m81_2/b[6] saout_m2_3v1024x8m81_2/b[7] saout_m2_3v1024x8m81_2/vss_uq4
+ saout_m2_3v1024x8m81_3/vdd saout_m2_3v1024x8m81_3/vdd_uq2 saout_m2_3v1024x8m81_3/vdd_uq1
+ pcb[5] saout_m2_3v1024x8m81_2/pcb_uq1 saout_m2_3v1024x8m81_2/bb[5] saout_m2_3v1024x8m81_2/mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/bb
+ saout_m2_3v1024x8m81_2/mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ saout_m2_3v1024x8m81_2/bb[2] GWE saout_m2_3v1024x8m81_2/bb[4] WEN[5] saout_m2_3v1024x8m81_2/bb[7]
+ saout_m2_3v1024x8m81_2/b[4] saout_m2_3v1024x8m81_3/men saout_R_m2_3v1024x8m81_3/vdd
+ saout_m2_3v1024x8m81_3/VDD saout_m2_3v1024x8m81_2/b[1] saout_m2_3v1024x8m81_2/bb[3]
+ saout_m2_3v1024x8m81_3/ypass[3] saout_m2_3v1024x8m81_3/ypass[6] saout_m2_3v1024x8m81_3/ypass[7]
+ saout_m2_3v1024x8m81_3/VDD_uq0 saout_m2_3v1024x8m81_3/ypass[5] saout_m2_3v1024x8m81_2/b[3]
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq0 saout_m2_3v1024x8m81_2/bb[6]
+ VSS saout_m2_3v1024x8m81
Xsaout_m2_3v1024x8m81_3 saout_m2_3v1024x8m81_3/ypass[1] saout_m2_3v1024x8m81_3/ypass[2]
+ saout_m2_3v1024x8m81_3/ypass[4] saout_m2_3v1024x8m81_3/ypass[0] saout_m2_3v1024x8m81_3/GWEN
+ d[4] q[4] saout_m2_3v1024x8m81_3/pcb saout_m2_3v1024x8m81_3/bb[0] saout_m2_3v1024x8m81_3/b[0]
+ saout_m2_3v1024x8m81_3/bb[1] saout_m2_3v1024x8m81_3/b[2] saout_m2_3v1024x8m81_3/b[5]
+ saout_m2_3v1024x8m81_3/b[6] saout_m2_3v1024x8m81_3/b[7] saout_m2_3v1024x8m81_3/vss_uq4
+ saout_m2_3v1024x8m81_3/vdd saout_m2_3v1024x8m81_3/vdd_uq2 saout_m2_3v1024x8m81_3/vdd_uq1
+ pcb[7] saout_m2_3v1024x8m81_3/pcb_uq1 saout_m2_3v1024x8m81_3/bb[5] saout_m2_3v1024x8m81_3/mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/bb
+ saout_m2_3v1024x8m81_3/mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ saout_m2_3v1024x8m81_3/bb[2] GWE saout_m2_3v1024x8m81_3/bb[4] WEN[7] saout_m2_3v1024x8m81_3/bb[7]
+ saout_m2_3v1024x8m81_3/b[4] saout_m2_3v1024x8m81_3/men saout_R_m2_3v1024x8m81_3/vdd
+ saout_m2_3v1024x8m81_3/VDD saout_m2_3v1024x8m81_3/b[1] saout_m2_3v1024x8m81_3/bb[3]
+ saout_m2_3v1024x8m81_3/ypass[3] saout_m2_3v1024x8m81_3/ypass[6] saout_m2_3v1024x8m81_3/ypass[7]
+ saout_m2_3v1024x8m81_3/VDD_uq0 saout_m2_3v1024x8m81_3/ypass[5] saout_m2_3v1024x8m81_3/b[3]
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq0 saout_m2_3v1024x8m81_3/bb[6]
+ VSS saout_m2_3v1024x8m81
Xrarray4_1024_3v1024x8m81_0 rarray4_1024_3v1024x8m81_0/m3_n1397_74227# WL[47] saout_m2_3v1024x8m81_2/bb[5]
+ rarray4_1024_3v1024x8m81_0/m3_n1397_64531# saout_m2_3v1024x8m81_3/b[2] saout_R_m2_3v1024x8m81_1/b[0]
+ saout_m2_3v1024x8m81_2/bb[6] saout_R_m2_3v1024x8m81_3/bb[2] saout_m2_3v1024x8m81_3/bb[4]
+ WL[4] saout_R_m2_3v1024x8m81_1/b[7] rarray4_1024_3v1024x8m81_0/m3_n1397_39793# rarray4_1024_3v1024x8m81_0/m3_n1397_41503#
+ saout_m2_3v1024x8m81_2/b[4] rarray4_1024_3v1024x8m81_0/m3_n1397_48775# saout_R_m2_3v1024x8m81_3/bb[7]
+ WL[3] rarray4_1024_3v1024x8m81_0/m3_n1397_61609# saout_m2_3v1024x8m81_2/mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/bb
+ WL[42] saout_m2_3v1024x8m81_3/bb[3] saout_m2_3v1024x8m81_2/b[1] saout_R_m2_3v1024x8m81_1/bb[4]
+ rarray4_1024_3v1024x8m81_0/m3_n1397_70591# rarray4_1024_3v1024x8m81_0/m3_n1397_26461#
+ saout_m2_3v1024x8m81_2/b[5] saout_m2_3v1024x8m81_3/bb[5] rarray4_1024_3v1024x8m81_0/m3_n1397_53125#
+ WL[28] rarray4_1024_3v1024x8m81_0/m3_n1397_51913# saout_R_m2_3v1024x8m81_3/b[5]
+ rarray4_1024_3v1024x8m81_0/m3_n1397_8779# saout_m2_3v1024x8m81_3/bb[2] rarray4_1024_3v1024x8m81_0/m3_n1397_22111#
+ WL[49] rarray4_1024_3v1024x8m81_0/m3_n1397_76153# rarray4_1024_3v1024x8m81_0/m3_n1397_40291#
+ saout_R_m2_3v1024x8m81_1/b[5] rarray4_1024_3v1024x8m81_0/m3_n1397_49987# WL[26]
+ WL[5] saout_R_m2_3v1024x8m81_3/b[2] rarray4_1024_3v1024x8m81_0/m3_n1397_47563# saout_R_m2_3v1024x8m81_3/bb[1]
+ WL[21] WL[32] WL[1] rarray4_1024_3v1024x8m81_0/m3_n1397_70093# rarray4_1024_3v1024x8m81_0/m3_n1397_57259#
+ saout_m2_3v1024x8m81_3/mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ saout_R_m2_3v1024x8m81_1/bb[7] saout_R_m2_3v1024x8m81_1/bb[2] rarray4_1024_3v1024x8m81_0/m3_n1397_62107#
+ saout_m2_3v1024x8m81_2/bb[3] saout_R_m2_3v1024x8m81_1/b[1] rarray4_1024_3v1024x8m81_0/m3_n1397_54337#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_19687# saout_R_m2_3v1024x8m81_1/b[6] WL[29]
+ rarray4_1024_3v1024x8m81_0/m3_n1397_71305# saout_m2_3v1024x8m81_3/b[6] saout_m2_3v1024x8m81_2/bb[4]
+ rarray4_1024_3v1024x8m81_0/m3_n1397_60895# rarray4_1024_3v1024x8m81_0/m3_n1397_48277#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_36655# rarray4_1024_3v1024x8m81_0/m3_n1397_59185#
+ WL[15] saout_R_m2_3v1024x8m81_3/bb[6] saout_m2_3v1024x8m81_2/bb[7] rarray4_1024_3v1024x8m81_0/m3_n1397_27673#
+ saout_m2_3v1024x8m81_3/b[3] saout_R_m2_3v1024x8m81_3/bb[4] rarray4_1024_3v1024x8m81_0/m3_n1397_57973#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_68881# rarray4_1024_3v1024x8m81_0/m3_n1397_13129#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_51199# saout_R_m2_3v1024x8m81_1/b[4] rarray4_1024_3v1024x8m81_0/m3_n1397_74941#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_35443# rarray4_1024_3v1024x8m81_0/m3_n1397_20899#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_43429# rarray4_1024_3v1024x8m81_0/m3_n1397_53623#
+ WL[19] saout_m2_3v1024x8m81_3/b[7] saout_R_m2_3v1024x8m81_1/bb[6] rarray4_1024_3v1024x8m81_0/m3_n1397_41005#
+ saout_m2_3v1024x8m81_3/b[5] rarray4_1024_3v1024x8m81_0/m3_n1397_73729# rarray4_1024_3v1024x8m81_0/m3_n1397_23323#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_77365# rarray4_1024_3v1024x8m81_0/m3_n1397_52411#
+ WL[59] WL[23] WL[24] saout_m2_3v1024x8m81_2/b[2] saout_R_m2_3v1024x8m81_3/b[0] saout_m2_3v1024x8m81_2/bb[2]
+ rarray4_1024_3v1024x8m81_0/m3_n1397_11917# WL[9] saout_m2_3v1024x8m81_2/mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ WL[54] rarray4_1024_3v1024x8m81_0/m3_n1397_69379# WL[22] WL[30] rarray4_1024_3v1024x8m81_0/m3_n1397_10705#
+ saout_R_m2_3v1024x8m81_3/bb[5] WL[7] rarray4_1024_3v1024x8m81_0/m3_n1397_67669#
+ saout_R_m2_3v1024x8m81_1/bb[3] WL[36] rarray4_1024_3v1024x8m81_0/m3_n1397_68167#
+ WL[61] WL[57] rarray4_1024_3v1024x8m81_0/m3_n1397_56047# WL[34] saout_R_m2_3v1024x8m81_1/bb[5]
+ saout_m2_3v1024x8m81_3/bb[1] saout_R_m2_3v1024x8m81_1/bb[0] rarray4_1024_3v1024x8m81_0/m3_n1397_73015#
+ WL[0] rarray4_1024_3v1024x8m81_0/m3_n1397_56761# WL[44] saout_m2_3v1024x8m81_3/b[1]
+ rarray4_1024_3v1024x8m81_0/m3_n1397_66955# WL[2] rarray4_1024_3v1024x8m81_0/m3_n1397_63319#
+ saout_R_m2_3v1024x8m81_3/bb[3] saout_m2_3v1024x8m81_3/bb[7] rarray4_1024_3v1024x8m81_0/m3_n1397_47065#
+ saout_m2_3v1024x8m81_3/b[4] rarray4_1024_3v1024x8m81_0/m3_n1397_24037# rarray4_1024_3v1024x8m81_0/m3_n1397_64033#
+ WL[46] rarray4_1024_3v1024x8m81_0/m3_n1397_46351# WL[55] rarray4_1024_3v1024x8m81_0/m3_n1397_72517#
+ saout_R_m2_3v1024x8m81_3/b[7] rarray4_1024_3v1024x8m81_0/m3_n1397_37867# saout_m2_3v1024x8m81_2/b[6]
+ rarray4_1024_3v1024x8m81_0/m3_n1397_50701# rarray4_1024_3v1024x8m81_0/m3_n1397_9493#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_54835# rarray4_1024_3v1024x8m81_0/m3_n1397_8281#
+ WL[27] WL[50] rarray4_1024_3v1024x8m81_0/m3_n1397_65743# rarray4_1024_3v1024x8m81_0/m3_n1397_71803#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_76651# saout_m2_3v1024x8m81_3/mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/bb
+ saout_R_m2_3v1024x8m81_3/b[3] saout_R_m2_3v1024x8m81_1/b[2] rarray4_1024_3v1024x8m81_0/m3_n1397_49489#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_5143# rarray4_1024_3v1024x8m81_0/m3_n1397_55549#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_28885# saout_m2_3v1024x8m81_2/b[3] rarray4_1024_3v1024x8m81_0/m3_n1397_59683#
+ saout_R_m2_3v1024x8m81_1/bb[1] rarray4_1024_3v1024x8m81_0/m3_n1397_6355# WL[52]
+ rarray4_1024_3v1024x8m81_0/m3_n1397_45853# rarray4_1024_3v1024x8m81_0/m3_n1397_62821#
+ WL[53] rarray4_1024_3v1024x8m81_0/m3_n1397_42715# saout_R_m2_3v1024x8m81_3/b[1]
+ saout_m2_3v1024x8m81_3/bb[6] saout_R_m2_3v1024x8m81_3/bb[0] saout_R_m2_3v1024x8m81_1/b[3]
+ rarray4_1024_3v1024x8m81_0/m3_n1397_44641# rarray4_1024_3v1024x8m81_0/m3_n1397_58471#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_45139# WL[11] rarray4_1024_3v1024x8m81_0/m3_n1397_39079#
+ WL[48] rarray4_1024_3v1024x8m81_0/m3_n1397_7567# saout_R_m2_3v1024x8m81_3/b[6] saout_m2_3v1024x8m81_2/b[7]
+ saout_m2_3v1024x8m81_2/bb[1] WL[25] rarray4_1024_3v1024x8m81_0/m3_n1397_25249# rarray4_1024_3v1024x8m81_0/m3_n1397_65245#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_3931# rarray4_1024_3v1024x8m81_0/m3_n1397_42217#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_43927# rarray4_1024_3v1024x8m81_0/m3_n1397_75439#
+ WL[40] WL[17] rarray4_1024_3v1024x8m81_0/m3_n1397_66457# rarray4_1024_3v1024x8m81_0/m3_n1397_24535#
+ WL[51] saout_m2_3v1024x8m81_3/vdd_uq3 saout_R_m2_3v1024x8m81_3/b[4] VSS rarray4_1024_3v1024x8m81_0/m3_n1397_60397#
+ rarray4_1024_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[0] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[1] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[2] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[3] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[4] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[5] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[6] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[7] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[8] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[9] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[10] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[11] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[12] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[13] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[14] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[15] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[16] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[17] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[18] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[19] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[20] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[21] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[22] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[23] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[24] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[25] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[26] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[27] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[28] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[29] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[30] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[31] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[32] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[33] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[34] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[35] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ dcap_103_novia_3v1024x8m81
Xrdummy_3v512x4_3v1024x8m81_0 VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS rarray4_1024_3v1024x8m81_0/m3_n1397_51199# saout_m2_3v1024x8m81_3/b[7] VSS rarray4_1024_3v1024x8m81_0/m3_n1397_77365#
+ WL[34] rarray4_1024_3v1024x8m81_0/m3_n1397_70591# saout_m2_3v1024x8m81_3/bb[7] saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3 WL[55] WL[26] rarray4_1024_3v1024x8m81_0/m3_n1397_43429#
+ VSS VSS VSS saout_R_m2_3v1024x8m81_3/b[7] tblhl saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_22111# saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/ypass[6] saout_R_m2_3v1024x8m81_3/bb[7] VSS WL[50] rarray4_1024_3v1024x8m81_0/m3_n1397_53125#
+ VSS rarray4_1024_3v1024x8m81_0/m3_n1397_49489# WL[50] VSS rarray4_1024_3v1024x8m81_0/m3_n1397_72517#
+ VSS VSS saout_m2_3v1024x8m81_2/b[7] saout_R_m2_3v1024x8m81_1/b[5] VSS saout_m2_3v1024x8m81_2/bb[2]
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_2/bb[7] saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_2/b[2] saout_R_m2_3v1024x8m81_1/bb[5] rarray4_1024_3v1024x8m81_0/m3_n1397_49987#
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_55549#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_26461# rarray4_1024_3v1024x8m81_0/m3_n1397_69379#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_25249# WL[9] VSS VSS VSS VSS saout_R_m2_3v1024x8m81_1/b[1]
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_R_m2_3v1024x8m81_3/b[1] WL[59] saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS saout_R_m2_3v1024x8m81_1/bb[1] saout_m2_3v1024x8m81_3/vdd_uq3 saout_R_m2_3v1024x8m81_3/bb[1]
+ saout_m2_3v1024x8m81_3/vdd saout_m2_3v1024x8m81_3/vdd_uq3 WL[0] saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS rarray4_1024_3v1024x8m81_0/m3_n1397_23323# WL[40] WL[23] VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS WL[46] saout_R_m2_3v1024x8m81_3/b[7] saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_51913#
+ VSS VSS rarray4_1024_3v1024x8m81_0/m3_n1397_71305# saout_R_m2_3v1024x8m81_3/bb[7]
+ saout_m2_3v1024x8m81_3/vdd_uq3 VSS rarray4_1024_3v1024x8m81_0/m3_n1397_45139# saout_m2_3v1024x8m81_3/vdd_uq3
+ WL[30] saout_m2_3v1024x8m81_3/vdd_uq3 VSS rarray4_1024_3v1024x8m81_0/m3_n1397_48775#
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_R_m2_3v1024x8m81_3/bb[0] saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_68167# saout_R_m2_3v1024x8m81_3/b[0] WL[36]
+ VSS VSS WL[51] rarray4_1024_3v1024x8m81_0/m3_n1397_51199# VSS WL[44] VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_2/b[3] saout_m2_3v1024x8m81_2/bb[6]
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_R_m2_3v1024x8m81_1/b[3]
+ saout_m2_3v1024x8m81_2/bb[3] saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_60895#
+ saout_m2_3v1024x8m81_2/b[6] saout_R_m2_3v1024x8m81_1/bb[3] rarray4_1024_3v1024x8m81_0/m3_n1397_50701#
+ WL[42] VSS saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_57259#
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 VSS WL[49] rarray4_1024_3v1024x8m81_0/m3_n1397_70093#
+ VSS rarray4_1024_3v1024x8m81_0/m3_n1397_8281# VSS VSS VSS saout_R_m2_3v1024x8m81_1/bb[4]
+ saout_R_m2_3v1024x8m81_3/bb[0] saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_R_m2_3v1024x8m81_1/b[4] rarray4_1024_3v1024x8m81_0/m3_n1397_66955#
+ tblhl saout_R_m2_3v1024x8m81_3/b[0] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_66955# saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_11917#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_24037# WL[19] saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3 VSS WL[47] saout_m2_3v1024x8m81_3/b[3]
+ VSS rarray4_1024_3v1024x8m81_0/m3_n1397_73015# saout_m2_3v1024x8m81_3/bb[3] VSS
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_44641# saout_m2_3v1024x8m81_3/vdd_uq3 WL[34]
+ VSS VSS rarray4_1024_3v1024x8m81_0/m3_n1397_49489# rarray4_1024_3v1024x8m81_0/m3_n1397_35443#
+ saout_R_m2_3v1024x8m81_3/bb[6] VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_68881# saout_R_m2_3v1024x8m81_3/b[6] VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_50701# WL[42]
+ VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_2/b[5] saout_m2_3v1024x8m81_2/mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/bb
+ saout_R_m2_3v1024x8m81_1/bb[2] rarray4_1024_3v1024x8m81_0/m3_n1397_65743# saout_m2_3v1024x8m81_2/bb[5]
+ saout_m2_3v1024x8m81_2/mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ saout_R_m2_3v1024x8m81_1/b[2] VSS rarray4_1024_3v1024x8m81_0/m3_n1397_60397# rarray4_1024_3v1024x8m81_0/m3_n1397_27673#
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 VSS rarray4_1024_3v1024x8m81_0/m3_n1397_56761#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_10705# WL[59] saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS VSS saout_R_m2_3v1024x8m81_1/bb[0] VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/bb
+ saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_66457# saout_m2_3v1024x8m81_3/mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ saout_R_m2_3v1024x8m81_1/b[0] saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_3931#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_37867# VSS VSS VSS rarray4_1024_3v1024x8m81_0/m3_n1397_40291#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_47563# rarray4_1024_3v1024x8m81_0/m3_n1397_67669#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_19687# WL[21] VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3 VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/b[5]
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/bb[5] rarray4_1024_3v1024x8m81_0/m3_n1397_72517#
+ saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_64531#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_46351# WL[36] VSS VSS WL[57] VSS saout_R_m2_3v1024x8m81_3/bb[4]
+ saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_R_m2_3v1024x8m81_3/b[4]
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_52411# saout_m2_3v1024x8m81_3/vdd_uq3 rdummy_3v512x4_3v1024x8m81_0/ypass_gate_3v1024x8m81_0_0/b
+ rarray4_1024_3v1024x8m81_0/m3_n1397_37867# VSS VSS WL[52] saout_m2_3v1024x8m81_2/bb[4]
+ saout_m2_3v1024x8m81_2/bb[4] VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_R_m2_3v1024x8m81_1/b[1]
+ rarray4_1024_3v1024x8m81_0/m3_n1397_46351# rarray4_1024_3v1024x8m81_0/m3_n1397_66457#
+ WL[0] saout_m2_3v1024x8m81_2/b[4] rarray4_1024_3v1024x8m81_0/m3_n1397_62107# VSS
+ VSS VSS saout_R_m2_3v1024x8m81_1/bb[1] saout_m2_3v1024x8m81_2/b[4] saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_58471# WL[53] WL[1] saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/b[1] saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_R_m2_3v1024x8m81_1/b[7] rarray4_1024_3v1024x8m81_0/m3_n1397_63319# saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_R_m2_3v1024x8m81_1/bb[7] VSS rarray4_1024_3v1024x8m81_0/m3_n1397_68167# saout_m2_3v1024x8m81_3/bb[1]
+ WL[61] rarray4_1024_3v1024x8m81_0/m3_n1397_5143# VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_48277#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_39793# WL[32] saout_m2_3v1024x8m81_3/vdd_uq3
+ WL[29] VSS VSS VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/bb[4]
+ saout_m2_3v1024x8m81_3/ypass[7] saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/b[4]
+ rarray4_1024_3v1024x8m81_0/m3_n1397_74227# WL[48] VSS VSS rarray4_1024_3v1024x8m81_0/m3_n1397_3931#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_45139# rarray4_1024_3v1024x8m81_0/m3_n1397_65245#
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_45853#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_13129# VSS VSS VSS VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_R_m2_3v1024x8m81_3/b[5] saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_R_m2_3v1024x8m81_3/bb[5]
+ saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_62107# saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_35443# saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq0
+ rarray4_1024_3v1024x8m81_0/m3_n1397_51913# VSS VSS WL[53] VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_2/bb[6] saout_m2_3v1024x8m81_2/b[3] VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_R_m2_3v1024x8m81_1/bb[0] saout_m2_3v1024x8m81_3/vdd_uq3 WL[1] rarray4_1024_3v1024x8m81_0/m3_n1397_47065#
+ saout_m2_3v1024x8m81_2/bb[3] saout_m2_3v1024x8m81_2/b[6] saout_R_m2_3v1024x8m81_1/b[0]
+ VSS VSS rarray4_1024_3v1024x8m81_0/m3_n1397_61609# saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS rarray4_1024_3v1024x8m81_0/m3_n1397_57973# saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_28885#
+ WL[44] VSS VSS saout_R_m2_3v1024x8m81_1/bb[2] VSS saout_m2_3v1024x8m81_3/bb[2] saout_m2_3v1024x8m81_3/vdd_uq3
+ WL[2] rarray4_1024_3v1024x8m81_0/m3_n1397_43927# rarray4_1024_3v1024x8m81_0/m3_n1397_64033#
+ saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_R_m2_3v1024x8m81_1/b[2] rarray4_1024_3v1024x8m81_0/m3_n1397_67669#
+ saout_m2_3v1024x8m81_3/b[2] VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/ypass[3]
+ VSS WL[4] VSS saout_m2_3v1024x8m81_3/vdd_uq2 rarray4_1024_3v1024x8m81_0/m3_n1397_41503#
+ WL[27] saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 VSS VSS saout_m2_3v1024x8m81_3/bb[6]
+ saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_60895# saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/b[6] rarray4_1024_3v1024x8m81_0/m3_n1397_73729#
+ WL[49] VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3 WL[7] rarray4_1024_3v1024x8m81_0/m3_n1397_45853#
+ saout_m2_3v1024x8m81_3/vdd_uq3 WL[24] VSS rarray4_1024_3v1024x8m81_0/m3_n1397_47563#
+ saout_m2_3v1024x8m81_3/vdd_uq3 VSS VSS VSS saout_R_m2_3v1024x8m81_3/b[3] saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_R_m2_3v1024x8m81_3/bb[3]
+ saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_42715# rarray4_1024_3v1024x8m81_0/m3_n1397_8779#
+ saout_m2_3v1024x8m81_3/ypass[4] rarray4_1024_3v1024x8m81_0/m3_n1397_62821# VSS rarray4_1024_3v1024x8m81_0/m3_n1397_53623#
+ VSS VSS WL[52] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS saout_m2_3v1024x8m81_2/b[7] saout_m2_3v1024x8m81_2/bb[2] saout_R_m2_3v1024x8m81_3/bb[6]
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_2/b[2]
+ saout_m2_3v1024x8m81_2/bb[7] saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_63319#
+ saout_R_m2_3v1024x8m81_3/b[6] VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 WL[61] rarray4_1024_3v1024x8m81_0/m3_n1397_59683#
+ saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_28885# VSS VSS
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/b[3]
+ rarray4_1024_3v1024x8m81_0/m3_n1397_44641# WL[3] saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 VSS VSS saout_m2_3v1024x8m81_3/bb[3] rarray4_1024_3v1024x8m81_0/m3_n1397_69379#
+ WL[2] VSS saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_41005#
+ VSS saout_m2_3v1024x8m81_3/b[7] rarray4_1024_3v1024x8m81_0/m3_n1397_41503# rarray4_1024_3v1024x8m81_0/m3_n1397_61609#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_6355# saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_75439#
+ saout_m2_3v1024x8m81_3/bb[7] VSS rarray4_1024_3v1024x8m81_0/m3_n1397_47065# saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 VSS VSS saout_R_m2_3v1024x8m81_3/bb[2] saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_R_m2_3v1024x8m81_3/b[2]
+ rdummy_3v512x4_3v1024x8m81_0/m2_16574_21# saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_9493# WL[21] rarray4_1024_3v1024x8m81_0/m3_n1397_43429#
+ VSS VSS rarray4_1024_3v1024x8m81_0/m3_n1397_53125# VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_R_m2_3v1024x8m81_1/b[5] saout_R_m2_3v1024x8m81_1/b[7] saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_R_m2_3v1024x8m81_3/bb[4] saout_m2_3v1024x8m81_3/ypass[0]
+ saout_R_m2_3v1024x8m81_1/bb[7] saout_R_m2_3v1024x8m81_1/bb[5] rarray4_1024_3v1024x8m81_0/m3_n1397_62821#
+ saout_R_m2_3v1024x8m81_3/b[4] saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS rarray4_1024_3v1024x8m81_0/m3_n1397_40291# WL[15] VSS VSS rarray4_1024_3v1024x8m81_0/m3_n1397_59185#
+ WL[5] rarray4_1024_3v1024x8m81_0/m3_n1397_59683# VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/b[5] saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/bb[5] rarray4_1024_3v1024x8m81_0/m3_n1397_68881#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_6355# VSS saout_m2_3v1024x8m81_3/vdd_uq3 VSS
+ saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_76651# rarray4_1024_3v1024x8m81_0/m3_n1397_24535#
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 VSS VSS WL[29] saout_m2_3v1024x8m81_3/b[1]
+ WL[11] saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_42217#
+ VSS VSS VSS saout_m2_3v1024x8m81_3/bb[1] rarray4_1024_3v1024x8m81_0/m3_n1397_74941#
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 WL[25] VSS rarray4_1024_3v1024x8m81_0/m3_n1397_39079#
+ saout_m2_3v1024x8m81_3/mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/bb rarray4_1024_3v1024x8m81_0/m3_n1397_5143#
+ saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_58471# saout_m2_3v1024x8m81_3/mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ saout_m2_3v1024x8m81_3/vdd_uq3 VSS WL[22] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ WL[28] VSS saout_m2_3v1024x8m81_3/vdd saout_R_m2_3v1024x8m81_3/b[5] saout_R_m2_3v1024x8m81_1/bb[6]
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_R_m2_3v1024x8m81_1/bb[6] saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_75439# saout_R_m2_3v1024x8m81_1/b[6] saout_R_m2_3v1024x8m81_1/b[6]
+ saout_R_m2_3v1024x8m81_3/bb[5] saout_m2_3v1024x8m81_3/vdd_uq3 VSS rarray4_1024_3v1024x8m81_0/m3_n1397_64531#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_41005# saout_m2_3v1024x8m81_3/vdd_uq3 VSS WL[25]
+ rarray4_1024_3v1024x8m81_0/m3_n1397_10705# saout_m2_3v1024x8m81_3/vdd_uq3 VSS VSS
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 WL[48] saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_60397#
+ WL[7] VSS VSS VSS saout_m2_3v1024x8m81_3/bb[4] saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_70591#
+ saout_m2_3v1024x8m81_3/b[4] WL[17] WL[4] WL[17] saout_m2_3v1024x8m81_3/vdd_uq3 VSS
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_57259# rarray4_1024_3v1024x8m81_0/m3_n1397_77365#
+ saout_m2_3v1024x8m81_3/vdd_uq3 WL[47] rarray4_1024_3v1024x8m81_0/m3_n1397_19687#
+ VSS VSS VSS VSS WL[30] rdummy_3v512x4_3v1024x8m81_0/ypass_gate_3v1024x8m81_0_0/b
+ saout_m2_3v1024x8m81_3/bb[2] saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/b[2]
+ rarray4_1024_3v1024x8m81_0/m3_n1397_76651# saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_74227# rarray4_1024_3v1024x8m81_0/m3_n1397_42715#
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 VSS rarray4_1024_3v1024x8m81_0/m3_n1397_24037#
+ saout_m2_3v1024x8m81_3/vdd_uq3 VSS VSS rarray4_1024_3v1024x8m81_0/m3_n1397_39793#
+ WL[23] WL[9] VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_2/b[5]
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_2/bb[5]
+ saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_59185# VSS rarray4_1024_3v1024x8m81_0/m3_n1397_48775#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_25249# VSS rarray4_1024_3v1024x8m81_0/m3_n1397_7567#
+ VSS WL[40] VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_R_m2_3v1024x8m81_3/b[3]
+ saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_56047#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_76153# VSS saout_R_m2_3v1024x8m81_3/bb[3] VSS
+ rarray4_1024_3v1024x8m81_0/m3_n1397_64033# WL[26] VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_54835# WL[46] WL[11] VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS saout_m2_3v1024x8m81_3/bb[6] saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_73015#
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_70093# WL[27]
+ saout_m2_3v1024x8m81_3/b[6] rarray4_1024_3v1024x8m81_0/m3_n1397_11917# VSS WL[5]
+ WL[15] VSS VSS VSS VSS rarray4_1024_3v1024x8m81_0/m3_n1397_57973# WL[55] saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_23323# VSS VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_R_m2_3v1024x8m81_3/b[1] rarray4_1024_3v1024x8m81_0/m3_n1397_76153# saout_R_m2_3v1024x8m81_3/bb[1]
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS rarray4_1024_3v1024x8m81_0/m3_n1397_54835# rarray4_1024_3v1024x8m81_0/m3_n1397_74941#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_42217# WL[32] VSS VSS VSS WL[24] VSS saout_m2_3v1024x8m81_2/b[1]
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_2/bb[1]
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/ypass[5] saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_48277# rarray4_1024_3v1024x8m81_0/m3_n1397_36655#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_26461# VSS WL[19] VSS rarray4_1024_3v1024x8m81_0/m3_n1397_8281#
+ saout_m2_3v1024x8m81_2/mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/bb VSS VSS
+ saout_R_m2_3v1024x8m81_1/b[3] VSS rarray4_1024_3v1024x8m81_0/m3_n1397_56761# saout_R_m2_3v1024x8m81_1/bb[3]
+ saout_m2_3v1024x8m81_2/mux821_3v1024x8m81_0/ypass_gate_a_3v1024x8m81_0/pmos_5p0431059130201_3v1024x8m81_0/D
+ rarray4_1024_3v1024x8m81_0/m3_n1397_65743# VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_54337# rarray4_1024_3v1024x8m81_0/m3_n1397_39079#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_9493# VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_53623# rarray4_1024_3v1024x8m81_0/m3_n1397_73729#
+ VSS VSS rarray4_1024_3v1024x8m81_0/m3_n1397_71803# saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 WL[28] rarray4_1024_3v1024x8m81_0/m3_n1397_8779#
+ VSS VSS VSS rarray4_1024_3v1024x8m81_0/m3_n1397_27673# rarray4_1024_3v1024x8m81_0/m3_n1397_22111#
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_20899#
+ VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 WL[54] rarray4_1024_3v1024x8m81_0/m3_n1397_55549#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_43927# rdummy_3v512x4_3v1024x8m81_0/ypass_gate_3v1024x8m81_0_0/pcb
+ WL[22] VSS VSS VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_52411#
+ VSS WL[54] rarray4_1024_3v1024x8m81_0/m3_n1397_49987# VSS rarray4_1024_3v1024x8m81_0/m3_n1397_13129#
+ rarray4_1024_3v1024x8m81_0/m3_n1397_71803# VSS saout_m2_3v1024x8m81_2/b[1] VSS VSS
+ saout_R_m2_3v1024x8m81_1/bb[4] saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/ypass[1]
+ saout_m2_3v1024x8m81_2/bb[1] rdummy_3v512x4_3v1024x8m81_0/m2_16574_77581# rarray4_1024_3v1024x8m81_0/m3_n1397_65245#
+ saout_R_m2_3v1024x8m81_1/b[4] VSS saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_56047#
+ saout_m2_3v1024x8m81_3/vdd_uq3 WL[57] WL[3] rarray4_1024_3v1024x8m81_0/m3_n1397_24535#
+ VSS VSS VSS VSS saout_R_m2_3v1024x8m81_3/bb[2] saout_m2_3v1024x8m81_3/vdd_uq3 saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_54337# saout_m2_3v1024x8m81_3/vdd_uq3 rarray4_1024_3v1024x8m81_0/m3_n1397_36655#
+ VSS VSS VSS saout_m2_3v1024x8m81_3/vdd_uq3 VSS saout_R_m2_3v1024x8m81_3/b[2] rarray4_1024_3v1024x8m81_0/m3_n1397_71305#
+ VSS rarray4_1024_3v1024x8m81_0/m3_n1397_7567# VSS VSS WL[51] saout_m2_3v1024x8m81_3/vdd_uq3
+ rarray4_1024_3v1024x8m81_0/m3_n1397_20899# saout_m2_3v1024x8m81_3/ypass[2] saout_m2_3v1024x8m81_3/vdd_uq3
+ rdummy_3v512x4_3v1024x8m81
Xsaout_R_m2_3v1024x8m81_1 saout_m2_3v1024x8m81_3/ypass[1] saout_m2_3v1024x8m81_3/ypass[4]
+ saout_m2_3v1024x8m81_3/ypass[5] saout_m2_3v1024x8m81_3/GWEN din[7] saout_R_m2_3v1024x8m81_1/b[0]
+ saout_R_m2_3v1024x8m81_1/bb[7] q[7] saout_R_m2_3v1024x8m81_1/vss_uq6 saout_m2_3v1024x8m81_3/vdd_uq1
+ saout_m2_3v1024x8m81_3/VDD saout_R_m2_3v1024x8m81_1/vdd_uq2 saout_R_m2_3v1024x8m81_1/vdd_uq4
+ saout_R_m2_3v1024x8m81_1/vdd_uq6 saout_R_m2_3v1024x8m81_1/b[1] saout_R_m2_3v1024x8m81_1/b[5]
+ saout_R_m2_3v1024x8m81_1/bb[6] saout_R_m2_3v1024x8m81_1/bb[2] saout_R_m2_3v1024x8m81_1/b[7]
+ saout_R_m2_3v1024x8m81_1/bb[5] GWE saout_m2_3v1024x8m81_3/ypass[7] saout_R_m2_3v1024x8m81_1/bb[3]
+ WEN[4] saout_R_m2_3v1024x8m81_1/bb[0] saout_R_m2_3v1024x8m81_1/b[3] pcb[4] saout_m2_3v1024x8m81_3/men
+ saout_R_m2_3v1024x8m81_3/vdd saout_m2_3v1024x8m81_3/VDD_uq0 saout_R_m2_3v1024x8m81_1/b[2]
+ saout_m2_3v1024x8m81_3/vdd_uq2 saout_m2_3v1024x8m81_3/vdd saout_R_m2_3v1024x8m81_1/b[6]
+ saout_R_m2_3v1024x8m81_1/bb[4] saout_m2_3v1024x8m81_3/ypass[3] saout_m2_3v1024x8m81_3/ypass[2]
+ saout_m2_3v1024x8m81_3/ypass[6] saout_m2_3v1024x8m81_3/ypass[0] saout_R_m2_3v1024x8m81_1/b[4]
+ saout_m2_3v1024x8m81_3/vdd_uq0 VSS saout_R_m2_3v1024x8m81_1/bb[1] saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_R_m2_3v1024x8m81
Xsaout_R_m2_3v1024x8m81_3 saout_m2_3v1024x8m81_3/ypass[1] saout_m2_3v1024x8m81_3/ypass[4]
+ saout_m2_3v1024x8m81_3/ypass[5] saout_m2_3v1024x8m81_3/GWEN din[5] saout_R_m2_3v1024x8m81_3/b[0]
+ saout_R_m2_3v1024x8m81_3/bb[7] q[5] saout_R_m2_3v1024x8m81_3/vss_uq6 saout_m2_3v1024x8m81_3/vdd_uq1
+ saout_m2_3v1024x8m81_3/VDD saout_R_m2_3v1024x8m81_3/vdd_uq2 saout_R_m2_3v1024x8m81_3/vdd_uq4
+ saout_R_m2_3v1024x8m81_3/vdd_uq6 saout_R_m2_3v1024x8m81_3/b[1] saout_R_m2_3v1024x8m81_3/b[5]
+ saout_R_m2_3v1024x8m81_3/bb[6] saout_R_m2_3v1024x8m81_3/bb[2] saout_R_m2_3v1024x8m81_3/b[7]
+ saout_R_m2_3v1024x8m81_3/bb[5] GWE saout_m2_3v1024x8m81_3/ypass[7] saout_R_m2_3v1024x8m81_3/bb[3]
+ WEN[6] saout_R_m2_3v1024x8m81_3/bb[0] saout_R_m2_3v1024x8m81_3/b[3] pcb[6] saout_m2_3v1024x8m81_3/men
+ saout_R_m2_3v1024x8m81_3/vdd saout_m2_3v1024x8m81_3/VDD_uq0 saout_R_m2_3v1024x8m81_3/b[2]
+ saout_m2_3v1024x8m81_3/vdd_uq2 saout_m2_3v1024x8m81_3/vdd saout_R_m2_3v1024x8m81_3/b[6]
+ saout_R_m2_3v1024x8m81_3/bb[4] saout_m2_3v1024x8m81_3/ypass[3] saout_m2_3v1024x8m81_3/ypass[2]
+ saout_m2_3v1024x8m81_3/ypass[6] saout_m2_3v1024x8m81_3/ypass[0] saout_R_m2_3v1024x8m81_3/b[4]
+ saout_m2_3v1024x8m81_3/vdd_uq0 VSS saout_R_m2_3v1024x8m81_3/bb[1] saout_m2_3v1024x8m81_3/vdd_uq3
+ saout_R_m2_3v1024x8m81
.ends

.subckt Cell_array8x8_3v1024x8m81 b[8] b[24] bb[0] bb[9] b[26] b[1] bb[18] bb[2] b[28]
+ bb[8] b[3] bb[20] bb[25] bb[24] b[9] bb[4] b[21] bb[27] b[25] b[10] b[5] bb[17]
+ bb[22] bb[29] bb[26] wl[63] b[11] bb[1] b[12] wl[0] bb[6] b[23] b[30] b[27] wl[87]
+ b[2] b[14] b[7] wl[64] wl[51] bb[19] wl[40] wl[61] bb[28] wl[26] wl[1] wl[70] wl[4]
+ b[13] bb[3] b[16] wl[67] b[20] wl[18] wl[39] b[17] wl[54] wl[60] wl[88] b[29] wl[28]
+ wl[23] wl[117] b[18] b[4] wl[17] wl[55] wl[93] wl[44] wl[56] wl[58] bb[10] wl[62]
+ bb[21] wl[101] b[19] wl[94] wl[2] wl[72] wl[5] wl[91] bb[11] wl[105] wl[68] wl[41]
+ wl[19] wl[57] b[15] wl[69] bb[5] wl[95] wl[8] wl[103] wl[46] bb[12] wl[106] b[22]
+ wl[74] wl[29] wl[80] wl[79] wl[73] wl[7] wl[122] wl[90] wl[32] wl[24] b[31] wl[118]
+ bb[13] wl[25] wl[10] wl[110] wl[119] bb[30] wl[45] wl[124] wl[53] wl[11] b[6] wl[97]
+ wl[3] wl[96] wl[123] wl[102] wl[115] wl[121] wl[82] wl[30] wl[14] bb[14] wl[89]
+ wl[31] bb[23] wl[92] bb[31] wl[59] wl[65] wl[75] wl[9] wl[27] wl[34] wl[77] wl[108]
+ wl[42] wl[107] wl[78] wl[12] bb[15] wl[109] wl[112] wl[37] wl[111] wl[47] wl[43]
+ wl[126] wl[81] wl[36] wl[98] wl[13] wl[100] wl[104] wl[22] wl[71] wl[113] wl[6]
+ bb[7] wl[38] wl[99] wl[66] wl[20] wl[50] wl[114] wl[86] wl[125] wl[16] wl[84] wl[48]
+ wl[120] wl[83] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] wl[116] wl[33] wl[52] bb[16] wl[76] wl[85] wl[15] wl[21] wl[49] b[0] wl[127]
+ VSUBS
X018SRAM_cell1_2x_3v1024x8m81_0[0|0] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[1|0] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[2|0] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[3|0] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[4|0] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[5|0] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[6|0] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[7|0] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[8|0] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[9|0] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[10|0] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[11|0] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[12|0] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[13|0] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[14|0] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[15|0] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[16|0] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[17|0] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[18|0] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[19|0] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[20|0] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[21|0] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[22|0] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[23|0] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[24|0] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[25|0] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[26|0] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[27|0] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[28|0] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[29|0] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[30|0] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[31|0] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[32|0] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[33|0] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[34|0] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[35|0] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[36|0] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[37|0] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[38|0] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[39|0] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[40|0] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[41|0] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[42|0] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[43|0] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[44|0] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[45|0] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[46|0] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[47|0] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[48|0] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[49|0] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[50|0] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[51|0] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[52|0] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[53|0] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[54|0] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[55|0] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[56|0] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[57|0] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[58|0] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[59|0] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[60|0] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[61|0] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[62|0] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[63|0] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[7] bb[7]
+ wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[0|1] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[1|1] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[2|1] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[3|1] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[4|1] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[5|1] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[6|1] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[7|1] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[8|1] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[9|1] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[10|1] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[11|1] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[12|1] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[13|1] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[14|1] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[15|1] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[16|1] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[17|1] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[18|1] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[19|1] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[20|1] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[21|1] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[22|1] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[23|1] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[24|1] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[25|1] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[26|1] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[27|1] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[28|1] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[29|1] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[30|1] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[31|1] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[32|1] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[33|1] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[34|1] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[35|1] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[36|1] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[37|1] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[38|1] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[39|1] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[40|1] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[41|1] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[42|1] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[43|1] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[44|1] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[45|1] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[46|1] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[47|1] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[48|1] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[49|1] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[50|1] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[51|1] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[52|1] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[53|1] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[54|1] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[55|1] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[56|1] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[57|1] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[58|1] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[59|1] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[60|1] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[61|1] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[62|1] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[63|1] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[6]
+ b[6] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[0|2] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[1|2] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[2|2] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[3|2] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[4|2] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[5|2] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[6|2] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[7|2] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[8|2] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[9|2] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[10|2] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[11|2] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[12|2] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[13|2] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[14|2] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[15|2] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[16|2] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[17|2] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[18|2] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[19|2] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[20|2] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[21|2] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[22|2] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[23|2] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[24|2] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[25|2] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[26|2] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[27|2] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[28|2] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[29|2] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[30|2] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[31|2] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[32|2] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[33|2] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[34|2] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[35|2] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[36|2] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[37|2] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[38|2] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[39|2] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[40|2] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[41|2] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[42|2] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[43|2] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[44|2] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[45|2] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[46|2] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[47|2] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[48|2] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[49|2] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[50|2] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[51|2] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[52|2] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[53|2] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[54|2] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[55|2] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[56|2] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[57|2] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[58|2] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[59|2] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[60|2] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[61|2] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[62|2] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[63|2] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[5] bb[5]
+ wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[0|3] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[1|3] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[2|3] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[3|3] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[4|3] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[5|3] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[6|3] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[7|3] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[8|3] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[9|3] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[10|3] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[11|3] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[12|3] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[13|3] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[14|3] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[15|3] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[16|3] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[17|3] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[18|3] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[19|3] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[20|3] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[21|3] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[22|3] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[23|3] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[24|3] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[25|3] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[26|3] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[27|3] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[28|3] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[29|3] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[30|3] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[31|3] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[32|3] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[33|3] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[34|3] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[35|3] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[36|3] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[37|3] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[38|3] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[39|3] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[40|3] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[41|3] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[42|3] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[43|3] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[44|3] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[45|3] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[46|3] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[47|3] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[48|3] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[49|3] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[50|3] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[51|3] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[52|3] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[53|3] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[54|3] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[55|3] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[56|3] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[57|3] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[58|3] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[59|3] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[60|3] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[61|3] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[62|3] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[63|3] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[4]
+ b[4] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[0|4] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[1|4] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[2|4] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[3|4] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[4|4] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[5|4] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[6|4] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[7|4] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[8|4] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[9|4] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[10|4] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[11|4] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[12|4] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[13|4] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[14|4] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[15|4] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[16|4] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[17|4] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[18|4] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[19|4] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[20|4] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[21|4] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[22|4] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[23|4] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[24|4] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[25|4] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[26|4] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[27|4] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[28|4] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[29|4] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[30|4] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[31|4] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[32|4] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[33|4] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[34|4] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[35|4] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[36|4] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[37|4] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[38|4] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[39|4] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[40|4] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[41|4] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[42|4] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[43|4] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[44|4] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[45|4] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[46|4] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[47|4] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[48|4] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[49|4] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[50|4] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[51|4] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[52|4] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[53|4] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[54|4] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[55|4] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[56|4] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[57|4] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[58|4] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[59|4] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[60|4] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[61|4] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[62|4] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[63|4] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[3] bb[3]
+ wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[0|5] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[1|5] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[2|5] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[3|5] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[4|5] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[5|5] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[6|5] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[7|5] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[8|5] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[9|5] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[10|5] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[11|5] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[12|5] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[13|5] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[14|5] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[15|5] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[16|5] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[17|5] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[18|5] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[19|5] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[20|5] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[21|5] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[22|5] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[23|5] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[24|5] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[25|5] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[26|5] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[27|5] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[28|5] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[29|5] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[30|5] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[31|5] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[32|5] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[33|5] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[34|5] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[35|5] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[36|5] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[37|5] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[38|5] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[39|5] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[40|5] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[41|5] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[42|5] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[43|5] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[44|5] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[45|5] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[46|5] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[47|5] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[48|5] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[49|5] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[50|5] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[51|5] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[52|5] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[53|5] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[54|5] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[55|5] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[56|5] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[57|5] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[58|5] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[59|5] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[60|5] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[61|5] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[62|5] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[63|5] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[2]
+ b[2] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[0|6] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[1|6] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[2|6] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[3|6] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[4|6] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[5|6] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[6|6] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[7|6] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[8|6] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[9|6] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[10|6] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[11|6] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[12|6] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[13|6] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[14|6] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[15|6] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[16|6] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[17|6] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[18|6] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[19|6] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[20|6] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[21|6] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[22|6] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[23|6] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[24|6] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[25|6] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[26|6] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[27|6] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[28|6] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[29|6] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[30|6] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[31|6] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[32|6] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[33|6] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[34|6] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[35|6] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[36|6] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[37|6] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[38|6] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[39|6] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[40|6] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[41|6] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[42|6] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[43|6] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[44|6] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[45|6] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[46|6] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[47|6] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[48|6] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[49|6] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[50|6] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[51|6] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[52|6] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[53|6] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[54|6] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[55|6] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[56|6] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[57|6] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[58|6] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[59|6] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[60|6] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[61|6] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[62|6] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[63|6] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[1] bb[1]
+ wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[0|7] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[1|7] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[2|7] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[3|7] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[4|7] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[5|7] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[6|7] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[7|7] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[8|7] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[9|7] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[10|7] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[11|7] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[12|7] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[13|7] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[14|7] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[15|7] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[16|7] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[17|7] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[18|7] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[19|7] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[20|7] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[21|7] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[22|7] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[23|7] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[24|7] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[25|7] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[26|7] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[27|7] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[28|7] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[29|7] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[30|7] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[31|7] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[32|7] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[33|7] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[34|7] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[35|7] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[36|7] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[37|7] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[38|7] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[39|7] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[40|7] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[41|7] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[42|7] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[43|7] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[44|7] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[45|7] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[46|7] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[47|7] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[48|7] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[49|7] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[50|7] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[51|7] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[52|7] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[53|7] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[54|7] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[55|7] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[56|7] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[57|7] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[58|7] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[59|7] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[60|7] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[61|7] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[62|7] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_0[63|7] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[0]
+ b[0] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[0|0] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[1|0] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[2|0] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[3|0] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[4|0] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[5|0] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[6|0] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[7|0] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[8|0] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[9|0] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[10|0] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[11|0] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[12|0] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[13|0] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[14|0] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[15|0] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[16|0] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[17|0] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[18|0] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[19|0] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[20|0] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[21|0] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[22|0] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[23|0] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[24|0] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[25|0] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[26|0] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[27|0] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[28|0] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[29|0] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[30|0] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[31|0] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[32|0] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[33|0] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[34|0] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[35|0] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[36|0] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[37|0] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[38|0] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[39|0] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[40|0] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[41|0] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[42|0] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[43|0] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[44|0] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[45|0] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[46|0] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[47|0] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[48|0] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[49|0] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[50|0] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[51|0] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[52|0] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[53|0] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[54|0] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[55|0] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[56|0] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[57|0] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[58|0] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[59|0] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[60|0] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[61|0] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[62|0] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[63|0] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[23]
+ bb[23] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[0|1] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[1|1] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[2|1] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[3|1] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[4|1] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[5|1] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[6|1] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[7|1] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[8|1] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[9|1] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[10|1] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[11|1] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[12|1] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[13|1] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[14|1] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[15|1] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[16|1] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[17|1] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[18|1] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[19|1] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[20|1] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[21|1] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[22|1] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[23|1] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[24|1] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[25|1] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[26|1] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[27|1] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[28|1] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[29|1] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[30|1] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[31|1] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[32|1] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[33|1] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[34|1] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[35|1] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[36|1] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[37|1] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[38|1] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[39|1] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[40|1] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[41|1] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[42|1] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[43|1] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[44|1] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[45|1] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[46|1] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[47|1] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[48|1] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[49|1] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[50|1] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[51|1] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[52|1] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[53|1] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[54|1] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[55|1] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[56|1] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[57|1] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[58|1] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[59|1] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[60|1] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[61|1] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[62|1] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[63|1] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[22]
+ b[22] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[0|2] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[1|2] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[2|2] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[3|2] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[4|2] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[5|2] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[6|2] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[7|2] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[8|2] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[9|2] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[10|2] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[11|2] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[12|2] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[13|2] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[14|2] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[15|2] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[16|2] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[17|2] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[18|2] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[19|2] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[20|2] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[21|2] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[22|2] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[23|2] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[24|2] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[25|2] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[26|2] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[27|2] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[28|2] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[29|2] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[30|2] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[31|2] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[32|2] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[33|2] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[34|2] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[35|2] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[36|2] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[37|2] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[38|2] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[39|2] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[40|2] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[41|2] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[42|2] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[43|2] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[44|2] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[45|2] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[46|2] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[47|2] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[48|2] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[49|2] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[50|2] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[51|2] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[52|2] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[53|2] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[54|2] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[55|2] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[56|2] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[57|2] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[58|2] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[59|2] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[60|2] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[61|2] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[62|2] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[63|2] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[21]
+ bb[21] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[0|3] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[1|3] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[2|3] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[3|3] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[4|3] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[5|3] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[6|3] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[7|3] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[8|3] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[9|3] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[10|3] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[11|3] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[12|3] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[13|3] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[14|3] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[15|3] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[16|3] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[17|3] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[18|3] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[19|3] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[20|3] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[21|3] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[22|3] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[23|3] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[24|3] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[25|3] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[26|3] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[27|3] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[28|3] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[29|3] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[30|3] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[31|3] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[32|3] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[33|3] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[34|3] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[35|3] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[36|3] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[37|3] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[38|3] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[39|3] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[40|3] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[41|3] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[42|3] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[43|3] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[44|3] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[45|3] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[46|3] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[47|3] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[48|3] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[49|3] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[50|3] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[51|3] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[52|3] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[53|3] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[54|3] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[55|3] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[56|3] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[57|3] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[58|3] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[59|3] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[60|3] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[61|3] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[62|3] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[63|3] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[20]
+ b[20] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[0|4] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[1|4] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[2|4] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[3|4] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[4|4] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[5|4] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[6|4] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[7|4] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[8|4] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[9|4] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[10|4] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[11|4] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[12|4] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[13|4] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[14|4] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[15|4] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[16|4] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[17|4] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[18|4] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[19|4] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[20|4] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[21|4] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[22|4] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[23|4] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[24|4] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[25|4] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[26|4] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[27|4] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[28|4] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[29|4] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[30|4] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[31|4] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[32|4] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[33|4] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[34|4] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[35|4] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[36|4] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[37|4] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[38|4] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[39|4] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[40|4] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[41|4] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[42|4] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[43|4] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[44|4] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[45|4] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[46|4] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[47|4] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[48|4] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[49|4] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[50|4] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[51|4] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[52|4] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[53|4] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[54|4] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[55|4] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[56|4] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[57|4] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[58|4] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[59|4] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[60|4] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[61|4] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[62|4] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[63|4] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[19]
+ bb[19] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[0|5] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[1|5] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[2|5] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[3|5] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[4|5] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[5|5] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[6|5] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[7|5] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[8|5] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[9|5] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[10|5] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[11|5] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[12|5] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[13|5] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[14|5] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[15|5] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[16|5] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[17|5] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[18|5] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[19|5] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[20|5] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[21|5] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[22|5] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[23|5] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[24|5] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[25|5] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[26|5] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[27|5] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[28|5] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[29|5] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[30|5] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[31|5] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[32|5] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[33|5] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[34|5] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[35|5] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[36|5] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[37|5] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[38|5] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[39|5] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[40|5] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[41|5] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[42|5] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[43|5] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[44|5] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[45|5] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[46|5] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[47|5] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[48|5] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[49|5] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[50|5] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[51|5] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[52|5] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[53|5] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[54|5] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[55|5] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[56|5] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[57|5] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[58|5] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[59|5] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[60|5] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[61|5] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[62|5] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[63|5] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[18]
+ b[18] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[0|6] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[1|6] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[2|6] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[3|6] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[4|6] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[5|6] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[6|6] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[7|6] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[8|6] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[9|6] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[10|6] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[11|6] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[12|6] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[13|6] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[14|6] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[15|6] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[16|6] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[17|6] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[18|6] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[19|6] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[20|6] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[21|6] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[22|6] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[23|6] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[24|6] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[25|6] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[26|6] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[27|6] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[28|6] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[29|6] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[30|6] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[31|6] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[32|6] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[33|6] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[34|6] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[35|6] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[36|6] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[37|6] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[38|6] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[39|6] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[40|6] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[41|6] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[42|6] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[43|6] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[44|6] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[45|6] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[46|6] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[47|6] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[48|6] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[49|6] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[50|6] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[51|6] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[52|6] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[53|6] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[54|6] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[55|6] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[56|6] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[57|6] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[58|6] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[59|6] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[60|6] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[61|6] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[62|6] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[63|6] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[17]
+ bb[17] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[0|7] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[1|7] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[2|7] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[3|7] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[4|7] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[5|7] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[6|7] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[7|7] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[8|7] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[9|7] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[10|7] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[11|7] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[12|7] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[13|7] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[14|7] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[15|7] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[16|7] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[17|7] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[18|7] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[19|7] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[20|7] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[21|7] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[22|7] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[23|7] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[24|7] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[25|7] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[26|7] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[27|7] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[28|7] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[29|7] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[30|7] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[31|7] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[32|7] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[33|7] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[34|7] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[35|7] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[36|7] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[37|7] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[38|7] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[39|7] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[40|7] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[41|7] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[42|7] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[43|7] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[44|7] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[45|7] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[46|7] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[47|7] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[48|7] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[49|7] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[50|7] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[51|7] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[52|7] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[53|7] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[54|7] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[55|7] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[56|7] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[57|7] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[58|7] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[59|7] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[60|7] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[61|7] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[62|7] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_1[63|7] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[16]
+ b[16] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[0|0] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[1|0] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[2|0] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[3|0] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[4|0] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[5|0] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[6|0] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[7|0] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[8|0] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[9|0] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[10|0] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[11|0] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[12|0] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[13|0] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[14|0] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[15|0] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[16|0] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[17|0] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[18|0] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[19|0] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[20|0] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[21|0] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[22|0] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[23|0] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[24|0] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[25|0] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[26|0] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[27|0] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[28|0] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[29|0] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[30|0] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[31|0] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[32|0] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[33|0] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[34|0] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[35|0] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[36|0] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[37|0] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[38|0] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[39|0] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[40|0] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[41|0] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[42|0] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[43|0] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[44|0] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[45|0] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[46|0] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[47|0] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[48|0] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[49|0] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[50|0] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[51|0] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[52|0] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[53|0] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[54|0] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[55|0] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[56|0] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[57|0] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[58|0] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[59|0] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[60|0] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[61|0] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[62|0] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[63|0] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[31]
+ b[31] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[0|1] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[1|1] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[2|1] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[3|1] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[4|1] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[5|1] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[6|1] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[7|1] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[8|1] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[9|1] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[10|1] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[11|1] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[12|1] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[13|1] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[14|1] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[15|1] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[16|1] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[17|1] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[18|1] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[19|1] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[20|1] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[21|1] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[22|1] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[23|1] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[24|1] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[25|1] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[26|1] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[27|1] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[28|1] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[29|1] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[30|1] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[31|1] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[32|1] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[33|1] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[34|1] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[35|1] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[36|1] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[37|1] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[38|1] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[39|1] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[40|1] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[41|1] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[42|1] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[43|1] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[44|1] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[45|1] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[46|1] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[47|1] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[48|1] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[49|1] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[50|1] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[51|1] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[52|1] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[53|1] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[54|1] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[55|1] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[56|1] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[57|1] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[58|1] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[59|1] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[60|1] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[61|1] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[62|1] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[63|1] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[30]
+ bb[30] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[0|2] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[1|2] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[2|2] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[3|2] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[4|2] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[5|2] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[6|2] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[7|2] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[8|2] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[9|2] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[10|2] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[11|2] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[12|2] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[13|2] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[14|2] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[15|2] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[16|2] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[17|2] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[18|2] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[19|2] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[20|2] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[21|2] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[22|2] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[23|2] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[24|2] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[25|2] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[26|2] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[27|2] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[28|2] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[29|2] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[30|2] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[31|2] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[32|2] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[33|2] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[34|2] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[35|2] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[36|2] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[37|2] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[38|2] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[39|2] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[40|2] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[41|2] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[42|2] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[43|2] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[44|2] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[45|2] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[46|2] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[47|2] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[48|2] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[49|2] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[50|2] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[51|2] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[52|2] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[53|2] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[54|2] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[55|2] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[56|2] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[57|2] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[58|2] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[59|2] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[60|2] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[61|2] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[62|2] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[63|2] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[29]
+ b[29] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[0|3] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[1|3] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[2|3] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[3|3] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[4|3] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[5|3] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[6|3] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[7|3] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[8|3] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[9|3] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[10|3] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[11|3] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[12|3] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[13|3] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[14|3] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[15|3] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[16|3] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[17|3] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[18|3] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[19|3] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[20|3] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[21|3] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[22|3] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[23|3] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[24|3] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[25|3] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[26|3] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[27|3] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[28|3] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[29|3] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[30|3] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[31|3] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[32|3] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[33|3] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[34|3] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[35|3] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[36|3] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[37|3] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[38|3] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[39|3] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[40|3] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[41|3] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[42|3] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[43|3] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[44|3] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[45|3] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[46|3] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[47|3] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[48|3] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[49|3] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[50|3] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[51|3] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[52|3] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[53|3] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[54|3] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[55|3] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[56|3] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[57|3] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[58|3] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[59|3] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[60|3] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[61|3] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[62|3] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[63|3] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[28]
+ bb[28] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[0|4] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[1|4] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[2|4] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[3|4] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[4|4] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[5|4] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[6|4] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[7|4] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[8|4] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[9|4] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[10|4] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[11|4] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[12|4] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[13|4] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[14|4] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[15|4] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[16|4] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[17|4] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[18|4] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[19|4] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[20|4] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[21|4] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[22|4] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[23|4] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[24|4] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[25|4] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[26|4] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[27|4] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[28|4] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[29|4] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[30|4] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[31|4] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[32|4] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[33|4] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[34|4] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[35|4] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[36|4] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[37|4] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[38|4] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[39|4] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[40|4] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[41|4] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[42|4] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[43|4] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[44|4] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[45|4] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[46|4] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[47|4] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[48|4] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[49|4] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[50|4] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[51|4] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[52|4] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[53|4] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[54|4] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[55|4] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[56|4] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[57|4] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[58|4] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[59|4] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[60|4] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[61|4] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[62|4] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[63|4] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[27]
+ b[27] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[0|5] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[1|5] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[2|5] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[3|5] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[4|5] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[5|5] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[6|5] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[7|5] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[8|5] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[9|5] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[10|5] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[11|5] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[12|5] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[13|5] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[14|5] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[15|5] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[16|5] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[17|5] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[18|5] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[19|5] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[20|5] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[21|5] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[22|5] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[23|5] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[24|5] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[25|5] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[26|5] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[27|5] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[28|5] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[29|5] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[30|5] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[31|5] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[32|5] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[33|5] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[34|5] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[35|5] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[36|5] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[37|5] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[38|5] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[39|5] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[40|5] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[41|5] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[42|5] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[43|5] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[44|5] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[45|5] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[46|5] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[47|5] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[48|5] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[49|5] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[50|5] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[51|5] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[52|5] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[53|5] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[54|5] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[55|5] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[56|5] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[57|5] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[58|5] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[59|5] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[60|5] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[61|5] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[62|5] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[63|5] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[26]
+ bb[26] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[0|6] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[1|6] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[2|6] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[3|6] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[4|6] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[5|6] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[6|6] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[7|6] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[8|6] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[9|6] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[10|6] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[11|6] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[12|6] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[13|6] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[14|6] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[15|6] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[16|6] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[17|6] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[18|6] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[19|6] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[20|6] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[21|6] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[22|6] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[23|6] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[24|6] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[25|6] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[26|6] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[27|6] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[28|6] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[29|6] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[30|6] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[31|6] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[32|6] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[33|6] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[34|6] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[35|6] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[36|6] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[37|6] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[38|6] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[39|6] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[40|6] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[41|6] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[42|6] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[43|6] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[44|6] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[45|6] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[46|6] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[47|6] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[48|6] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[49|6] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[50|6] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[51|6] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[52|6] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[53|6] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[54|6] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[55|6] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[56|6] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[57|6] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[58|6] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[59|6] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[60|6] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[61|6] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[62|6] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[63|6] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[25]
+ b[25] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[0|7] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[1|7] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[2|7] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[3|7] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[4|7] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[5|7] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[6|7] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[7|7] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[8|7] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[9|7] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[10|7] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[11|7] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[12|7] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[13|7] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[14|7] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[15|7] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[16|7] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[17|7] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[18|7] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[19|7] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[20|7] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[21|7] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[22|7] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[23|7] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[24|7] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[25|7] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[26|7] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[27|7] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[28|7] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[29|7] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[30|7] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[31|7] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[32|7] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[33|7] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[34|7] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[35|7] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[36|7] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[37|7] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[38|7] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[39|7] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[40|7] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[41|7] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[42|7] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[43|7] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[44|7] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[45|7] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[46|7] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[47|7] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[48|7] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[49|7] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[50|7] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[51|7] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[52|7] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[53|7] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[54|7] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[55|7] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[56|7] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[57|7] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[58|7] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[59|7] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[60|7] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[61|7] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[62|7] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_2[63|7] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[24]
+ bb[24] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[0|0] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[1|0] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[2|0] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[3|0] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[4|0] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[5|0] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[6|0] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[7|0] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[8|0] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[9|0] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[10|0] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[11|0] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[12|0] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[13|0] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[14|0] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[15|0] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[16|0] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[17|0] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[18|0] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[19|0] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[20|0] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[21|0] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[22|0] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[23|0] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[24|0] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[25|0] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[26|0] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[27|0] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[28|0] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[29|0] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[30|0] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[31|0] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[32|0] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[33|0] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[34|0] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[35|0] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[36|0] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[37|0] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[38|0] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[39|0] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[40|0] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[41|0] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[42|0] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[43|0] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[44|0] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[45|0] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[46|0] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[47|0] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[48|0] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[49|0] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[50|0] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[51|0] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[52|0] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[53|0] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[54|0] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[55|0] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[56|0] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[57|0] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[58|0] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[59|0] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[60|0] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[61|0] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[62|0] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[63|0] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[15]
+ b[15] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[0|1] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[1|1] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[2|1] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[3|1] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[4|1] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[5|1] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[6|1] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[7|1] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[8|1] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[9|1] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[10|1] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[11|1] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[12|1] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[13|1] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[14|1] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[15|1] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[16|1] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[17|1] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[18|1] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[19|1] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[20|1] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[21|1] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[22|1] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[23|1] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[24|1] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[25|1] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[26|1] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[27|1] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[28|1] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[29|1] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[30|1] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[31|1] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[32|1] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[33|1] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[34|1] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[35|1] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[36|1] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[37|1] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[38|1] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[39|1] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[40|1] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[41|1] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[42|1] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[43|1] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[44|1] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[45|1] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[46|1] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[47|1] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[48|1] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[49|1] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[50|1] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[51|1] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[52|1] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[53|1] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[54|1] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[55|1] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[56|1] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[57|1] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[58|1] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[59|1] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[60|1] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[61|1] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[62|1] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[63|1] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[14]
+ bb[14] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[0|2] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[1|2] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[2|2] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[3|2] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[4|2] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[5|2] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[6|2] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[7|2] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[8|2] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[9|2] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[10|2] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[11|2] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[12|2] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[13|2] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[14|2] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[15|2] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[16|2] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[17|2] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[18|2] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[19|2] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[20|2] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[21|2] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[22|2] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[23|2] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[24|2] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[25|2] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[26|2] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[27|2] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[28|2] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[29|2] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[30|2] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[31|2] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[32|2] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[33|2] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[34|2] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[35|2] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[36|2] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[37|2] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[38|2] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[39|2] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[40|2] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[41|2] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[42|2] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[43|2] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[44|2] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[45|2] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[46|2] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[47|2] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[48|2] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[49|2] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[50|2] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[51|2] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[52|2] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[53|2] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[54|2] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[55|2] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[56|2] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[57|2] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[58|2] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[59|2] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[60|2] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[61|2] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[62|2] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[63|2] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[13]
+ b[13] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[0|3] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[1|3] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[2|3] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[3|3] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[4|3] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[5|3] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[6|3] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[7|3] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[8|3] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[9|3] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[10|3] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[11|3] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[12|3] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[13|3] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[14|3] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[15|3] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[16|3] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[17|3] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[18|3] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[19|3] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[20|3] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[21|3] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[22|3] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[23|3] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[24|3] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[25|3] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[26|3] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[27|3] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[28|3] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[29|3] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[30|3] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[31|3] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[32|3] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[33|3] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[34|3] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[35|3] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[36|3] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[37|3] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[38|3] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[39|3] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[40|3] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[41|3] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[42|3] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[43|3] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[44|3] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[45|3] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[46|3] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[47|3] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[48|3] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[49|3] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[50|3] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[51|3] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[52|3] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[53|3] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[54|3] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[55|3] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[56|3] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[57|3] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[58|3] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[59|3] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[60|3] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[61|3] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[62|3] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[63|3] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[12]
+ bb[12] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[0|4] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[1|4] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[2|4] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[3|4] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[4|4] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[5|4] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[6|4] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[7|4] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[8|4] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[9|4] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[10|4] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[11|4] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[12|4] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[13|4] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[14|4] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[15|4] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[16|4] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[17|4] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[18|4] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[19|4] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[20|4] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[21|4] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[22|4] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[23|4] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[24|4] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[25|4] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[26|4] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[27|4] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[28|4] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[29|4] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[30|4] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[31|4] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[32|4] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[33|4] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[34|4] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[35|4] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[36|4] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[37|4] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[38|4] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[39|4] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[40|4] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[41|4] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[42|4] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[43|4] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[44|4] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[45|4] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[46|4] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[47|4] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[48|4] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[49|4] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[50|4] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[51|4] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[52|4] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[53|4] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[54|4] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[55|4] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[56|4] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[57|4] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[58|4] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[59|4] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[60|4] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[61|4] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[62|4] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[63|4] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[11]
+ b[11] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[0|5] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[1|5] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[2|5] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[3|5] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[4|5] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[5|5] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[6|5] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[7|5] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[8|5] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[9|5] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[10|5] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[11|5] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[12|5] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[13|5] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[14|5] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[15|5] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[16|5] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[17|5] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[18|5] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[19|5] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[20|5] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[21|5] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[22|5] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[23|5] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[24|5] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[25|5] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[26|5] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[27|5] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[28|5] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[29|5] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[30|5] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[31|5] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[32|5] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[33|5] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[34|5] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[35|5] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[36|5] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[37|5] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[38|5] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[39|5] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[40|5] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[41|5] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[42|5] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[43|5] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[44|5] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[45|5] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[46|5] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[47|5] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[48|5] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[49|5] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[50|5] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[51|5] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[52|5] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[53|5] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[54|5] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[55|5] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[56|5] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[57|5] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[58|5] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[59|5] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[60|5] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[61|5] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[62|5] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[63|5] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[10]
+ bb[10] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[0|6] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[1|6] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[2|6] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[3|6] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[4|6] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[5|6] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[6|6] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[7|6] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[8|6] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[9|6] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[10|6] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[11|6] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[12|6] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[13|6] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[14|6] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[15|6] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[16|6] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[17|6] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[18|6] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[19|6] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[20|6] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[21|6] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[22|6] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[23|6] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[24|6] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[25|6] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[26|6] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[27|6] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[28|6] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[29|6] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[30|6] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[31|6] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[32|6] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[33|6] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[34|6] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[35|6] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[36|6] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[37|6] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[38|6] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[39|6] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[40|6] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[41|6] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[42|6] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[43|6] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[44|6] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[45|6] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[46|6] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[47|6] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[48|6] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[49|6] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[50|6] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[51|6] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[52|6] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[53|6] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[54|6] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[55|6] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[56|6] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[57|6] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[58|6] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[59|6] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[60|6] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[61|6] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[62|6] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[63|6] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# bb[9]
+ b[9] wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[0|7] wl[0] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[1]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[0] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[1] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[1|7] wl[2] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[3]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[2] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[3] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[2|7] wl[4] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[5]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[4] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[5] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[3|7] wl[6] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[7]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[6] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[7] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[4|7] wl[8] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[9]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[8] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[9] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[5|7] wl[10] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[11]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[10] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[11] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[6|7] wl[12] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[13]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[12] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[13] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[7|7] wl[14] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[15]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[14] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[15] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[8|7] wl[16] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[17]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[16] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[17] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[9|7] wl[18] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[19]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[18] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[19] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[10|7] wl[20] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[21]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[20] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[21] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[11|7] wl[22] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[23]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[22] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[23] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[12|7] wl[24] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[25]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[24] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[25] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[13|7] wl[26] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[27]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[26] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[27] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[14|7] wl[28] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[29]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[28] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[29] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[15|7] wl[30] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[31]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[30] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[31] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[16|7] wl[32] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[33]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[32] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[33] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[17|7] wl[34] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[35]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[34] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[35] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[18|7] wl[36] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[37]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[36] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[37] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[19|7] wl[38] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[39]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[38] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[39] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[20|7] wl[40] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[41]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[40] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[41] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[21|7] wl[42] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[43]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[42] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[43] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[22|7] wl[44] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[45]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[44] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[45] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[23|7] wl[46] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[47]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[46] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[47] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[24|7] wl[48] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[49]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[48] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[49] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[25|7] wl[50] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[51]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[50] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[51] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[26|7] wl[52] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[53]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[52] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[53] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[27|7] wl[54] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[55]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[54] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[55] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[28|7] wl[56] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[57]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[56] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[57] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[29|7] wl[58] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[59]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[58] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[59] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[30|7] wl[60] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[61]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[60] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[61] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[31|7] wl[62] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[63]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[62] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[63] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[32|7] wl[64] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[65]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[64] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[65] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[33|7] wl[66] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[67]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[66] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[67] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[34|7] wl[68] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[69]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[68] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[69] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[35|7] wl[70] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[71]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[70] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[71] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[36|7] wl[72] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[73]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[72] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[73] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[37|7] wl[74] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[75]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[74] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[75] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[38|7] wl[76] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[77]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[76] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[77] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[39|7] wl[78] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[79]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[78] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[79] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[40|7] wl[80] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[81]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[80] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[81] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[41|7] wl[82] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[83]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[82] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[83] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[42|7] wl[84] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[85]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[84] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[85] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[43|7] wl[86] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[87]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[86] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[87] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[44|7] wl[88] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[89]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[88] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[89] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[45|7] wl[90] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[91]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[90] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[91] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[46|7] wl[92] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[93]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[92] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[93] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[47|7] wl[94] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[95]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[94] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[95] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[48|7] wl[96] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[97]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[96] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[97] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[49|7] wl[98] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[99]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[98] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[99] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[50|7] wl[100] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[101]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[100] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[101] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[51|7] wl[102] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[103]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[102] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[103] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[52|7] wl[104] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[105]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[104] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[105] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[53|7] wl[106] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[107]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[106] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[107] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[54|7] wl[108] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[109]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[108] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[109] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[55|7] wl[110] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[111]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[110] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[111] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[56|7] wl[112] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[113]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[112] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[113] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[57|7] wl[114] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[115]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[114] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[115] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[58|7] wl[116] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[117]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[116] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[117] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[59|7] wl[118] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[119]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[118] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[119] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[60|7] wl[120] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[121]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[120] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[121] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[61|7] wl[122] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[123]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[122] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[123] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[62|7] wl[124] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[125]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[124] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[125] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
X018SRAM_cell1_2x_3v1024x8m81_3[63|7] wl[126] 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# wl[127]
+ 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512# b[8] bb[8]
+ wl[126] VSUBS 018SRAM_strap1_2x_3v1024x8m81_3[9]/018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ wl[127] VSUBS VSUBS x018SRAM_cell1_2x_3v1024x8m81
.ends

.subckt col_1024a_3v1024x8m81 WL[3] ypass[0] ypass[1] ypass[3] ypass[4] ypass[5] VDD
+ WL[32] WL[31] WL[30] WL[23] WL[22] WL[57] WL[20] WL[48] WL[12] WL[11] WL[50] WL[51]
+ WL[41] WL[40] WL[10] WL[43] WL[35] WL[34] WL[37] WL[33] WL[38] WL[36] WL[5] WL[18]
+ WL[55] WL[53] WL[17] WL[54] WL[52] WL[127] WL[61] WL[15] WL[14] WL[13] WL[0] ypass[2]
+ WL[25] b[16] b[19] din[1] din[3] din[2] din[0] q[0] q[1] q[2] q[3] b[17] b[14] b[8]
+ bb[8] bb[10] bb[11] bb[12] bb[13] bb[14] bb[15] bb[16] bb[24] bb[25] bb[27] bb[29]
+ bb[30] bb[31] b[30] b[24] b[0] b[18] pcb[0] pcb[1] pcb[3] pcb[2] WEN[3] WEN[2] WEN[0]
+ VDD_uq5 Cell_array8x8_3v1024x8m81_0/wl[81] WL[39] Cell_array8x8_3v1024x8m81_0/wl[108]
+ Cell_array8x8_3v1024x8m81_0/wl[126] Cell_array8x8_3v1024x8m81_0/wl[75] Cell_array8x8_3v1024x8m81_0/wl[93]
+ Cell_array8x8_3v1024x8m81_0/wl[111] Cell_array8x8_3v1024x8m81_0/wl[70] Cell_array8x8_3v1024x8m81_0/b[8]
+ Cell_array8x8_3v1024x8m81_0/wl[88] Cell_array8x8_3v1024x8m81_0/wl[90] Cell_array8x8_3v1024x8m81_0/wl[124]
+ Cell_array8x8_3v1024x8m81_0/wl[73] Cell_array8x8_3v1024x8m81_0/wl[91] Cell_array8x8_3v1024x8m81_0/wl[118]
+ Cell_array8x8_3v1024x8m81_0/wl[109] ypass[6] Cell_array8x8_3v1024x8m81_0/wl[68]
+ ypass[7] Cell_array8x8_3v1024x8m81_0/wl[86] Cell_array8x8_3v1024x8m81_0/wl[104]
+ m3_n771_22409# men Cell_array8x8_3v1024x8m81_0/wl[71] Cell_array8x8_3v1024x8m81_0/wl[98]
+ WL[1] bb[0] Cell_array8x8_3v1024x8m81_0/wl[89] Cell_array8x8_3v1024x8m81_0/wl[116]
+ WL[21] Cell_array8x8_3v1024x8m81_0/wl[106] Cell_array8x8_3v1024x8m81_0/wl[107] saout_R_m2_3v1024x8m81_0/vdd_uq4
+ bb[20] Cell_array8x8_3v1024x8m81_0/wl[66] Cell_array8x8_3v1024x8m81_0/wl[125] bb[2]
+ Cell_array8x8_3v1024x8m81_0/bb[24] Cell_array8x8_3v1024x8m81_0/wl[84] b[9] Cell_array8x8_3v1024x8m81_0/wl[102]
+ b[21] Cell_array8x8_3v1024x8m81_0/wl[119] bb[4] Cell_array8x8_3v1024x8m81_0/wl[78]
+ Cell_array8x8_3v1024x8m81_0/wl[120] WL[8] b[5] Cell_array8x8_3v1024x8m81_0/wl[96]
+ WL[28] bb[22] Cell_array8x8_3v1024x8m81_0/wl[87] Cell_array8x8_3v1024x8m81_0/wl[114]
+ bb[26] Cell_array8x8_3v1024x8m81_0/b[24] WL[46] Cell_array8x8_3v1024x8m81_0/wl[105]
+ bb[1] bb[6] Cell_array8x8_3v1024x8m81_0/wl[64] b[25] Cell_array8x8_3v1024x8m81_0/wl[123]
+ b[23] Cell_array8x8_3v1024x8m81_0/bb[8] Cell_array8x8_3v1024x8m81_0/wl[82] b[26]
+ b[7] bb[9] WL[58] Cell_array8x8_3v1024x8m81_0/wl[100] Cell_array8x8_3v1024x8m81_0/wl[117]
+ b[27] WL[49] Cell_array8x8_3v1024x8m81_0/wl[122] Cell_array8x8_3v1024x8m81_0/wl[76]
+ bb[28] WL[6] b[28] Cell_array8x8_3v1024x8m81_0/wl[67] b[13] Cell_array8x8_3v1024x8m81_0/wl[94]
+ bb[3] WL[26] VDD_uq2 Cell_array8x8_3v1024x8m81_0/wl[85] b[20] Cell_array8x8_3v1024x8m81_0/wl[112]
+ WL[44] b[29] Cell_array8x8_3v1024x8m81_0/wl[103] WL[62] Cell_array8x8_3v1024x8m81_0/wl[121]
+ Cell_array8x8_3v1024x8m81_0/wl[79] bb[17] WL[9] bb[21] Cell_array8x8_3v1024x8m81_0/wl[80]
+ VDD_uq4 Cell_array8x8_3v1024x8m81_0/wl[97] bb[18] WL[29] WL[56] Cell_array8x8_3v1024x8m81_0/wl[115]
+ b[15] bb[5] saout_m2_3v1024x8m81_4/GWEN WL[47] bb[19] Cell_array8x8_3v1024x8m81_0/wl[74]
+ b[22] WL[4] VDD_uq1 Cell_array8x8_3v1024x8m81_0/wl[65] b[31] Cell_array8x8_3v1024x8m81_0/wl[92]
+ GWE Cell_array8x8_3v1024x8m81_0/wl[99] VDD_uq0 WL[24] WEN[1] b[6] Cell_array8x8_3v1024x8m81_0/wl[110]
+ WL[42] bb[23] VDD_uq3 Cell_array8x8_3v1024x8m81_0/wl[101] WL[59] Cell_array8x8_3v1024x8m81_0/wl[83]
+ WL[60] WL[16] Cell_array8x8_3v1024x8m81_0/wl[77] b[1] b[10] Cell_array8x8_3v1024x8m81_0/wl[69]
+ bb[7] WL[7] Cell_array8x8_3v1024x8m81_0/wl[95] b[2] b[11] WL[27] Cell_array8x8_3v1024x8m81_0/wl[113]
+ b[3] b[12] WL[45] Cell_array8x8_3v1024x8m81_0/wl[72] WL[2] VDD_uq6 WL[19] Cell_array8x8_3v1024x8m81_0/wl[63]
+ VSS b[4]
Xsaout_m2_3v1024x8m81_3 ypass[1] ypass[2] ypass[4] ypass[0] saout_m2_3v1024x8m81_4/GWEN
+ din[0] q[0] saout_m2_3v1024x8m81_3/pcb bb[24] b[24] bb[25] b[26] b[29] b[30] b[31]
+ saout_m2_3v1024x8m81_3/vss_uq4 VDD_uq3 VDD_uq4 VDD_uq2 saout_m2_3v1024x8m81_3/pcb_uq0
+ saout_m2_3v1024x8m81_3/pcb_uq1 bb[29] Cell_array8x8_3v1024x8m81_0/bb[24] Cell_array8x8_3v1024x8m81_0/b[24]
+ bb[26] GWE bb[28] WEN[3] bb[31] b[28] men VDD VDD_uq0 b[25] bb[27] ypass[3] ypass[6]
+ ypass[7] VDD_uq1 ypass[5] b[27] VDD_uq6 VDD_uq5 bb[30] VSS saout_m2_3v1024x8m81
Xsaout_m2_3v1024x8m81_4 ypass[1] ypass[2] ypass[4] ypass[0] saout_m2_3v1024x8m81_4/GWEN
+ din[2] q[2] saout_m2_3v1024x8m81_4/pcb bb[8] b[8] bb[9] b[10] b[13] b[14] b[15]
+ saout_m2_3v1024x8m81_4/vss_uq4 VDD_uq3 VDD_uq4 VDD_uq2 saout_m2_3v1024x8m81_4/pcb_uq0
+ saout_m2_3v1024x8m81_4/pcb_uq1 bb[13] Cell_array8x8_3v1024x8m81_0/bb[8] Cell_array8x8_3v1024x8m81_0/b[8]
+ bb[10] GWE bb[12] WEN[1] bb[15] b[12] men VDD VDD_uq0 b[9] bb[11] ypass[3] ypass[6]
+ ypass[7] VDD_uq1 ypass[5] b[11] VDD_uq6 VDD_uq5 bb[14] VSS saout_m2_3v1024x8m81
XCell_array8x8_3v1024x8m81_0 Cell_array8x8_3v1024x8m81_0/b[8] Cell_array8x8_3v1024x8m81_0/b[24]
+ bb[0] bb[9] b[26] b[1] bb[18] bb[2] b[28] Cell_array8x8_3v1024x8m81_0/bb[8] b[3]
+ bb[20] bb[25] Cell_array8x8_3v1024x8m81_0/bb[24] b[9] bb[4] b[21] bb[27] b[25] b[10]
+ b[5] bb[17] bb[22] bb[29] bb[26] Cell_array8x8_3v1024x8m81_0/wl[63] b[11] bb[1]
+ b[12] WL[0] bb[6] b[23] b[30] b[27] Cell_array8x8_3v1024x8m81_0/wl[87] b[2] b[14]
+ b[7] Cell_array8x8_3v1024x8m81_0/wl[64] WL[51] bb[19] WL[40] WL[61] bb[28] WL[26]
+ WL[1] Cell_array8x8_3v1024x8m81_0/wl[70] WL[4] b[13] bb[3] b[16] Cell_array8x8_3v1024x8m81_0/wl[67]
+ b[20] WL[18] WL[39] b[17] WL[54] WL[60] Cell_array8x8_3v1024x8m81_0/wl[88] b[29]
+ WL[28] WL[23] Cell_array8x8_3v1024x8m81_0/wl[117] b[18] b[4] WL[17] WL[55] Cell_array8x8_3v1024x8m81_0/wl[93]
+ WL[44] WL[56] WL[58] bb[10] WL[62] bb[21] Cell_array8x8_3v1024x8m81_0/wl[101] b[19]
+ Cell_array8x8_3v1024x8m81_0/wl[94] WL[2] Cell_array8x8_3v1024x8m81_0/wl[72] WL[5]
+ Cell_array8x8_3v1024x8m81_0/wl[91] bb[11] Cell_array8x8_3v1024x8m81_0/wl[105] Cell_array8x8_3v1024x8m81_0/wl[68]
+ WL[41] WL[19] WL[57] b[15] Cell_array8x8_3v1024x8m81_0/wl[69] bb[5] Cell_array8x8_3v1024x8m81_0/wl[95]
+ WL[8] Cell_array8x8_3v1024x8m81_0/wl[103] WL[46] bb[12] Cell_array8x8_3v1024x8m81_0/wl[106]
+ b[22] Cell_array8x8_3v1024x8m81_0/wl[74] WL[29] Cell_array8x8_3v1024x8m81_0/wl[80]
+ Cell_array8x8_3v1024x8m81_0/wl[79] Cell_array8x8_3v1024x8m81_0/wl[73] WL[7] Cell_array8x8_3v1024x8m81_0/wl[122]
+ Cell_array8x8_3v1024x8m81_0/wl[90] WL[32] WL[24] b[31] Cell_array8x8_3v1024x8m81_0/wl[118]
+ bb[13] WL[25] WL[10] Cell_array8x8_3v1024x8m81_0/wl[110] Cell_array8x8_3v1024x8m81_0/wl[119]
+ bb[30] WL[45] Cell_array8x8_3v1024x8m81_0/wl[124] WL[53] WL[11] b[6] Cell_array8x8_3v1024x8m81_0/wl[97]
+ WL[3] Cell_array8x8_3v1024x8m81_0/wl[96] Cell_array8x8_3v1024x8m81_0/wl[123] Cell_array8x8_3v1024x8m81_0/wl[102]
+ Cell_array8x8_3v1024x8m81_0/wl[115] Cell_array8x8_3v1024x8m81_0/wl[121] Cell_array8x8_3v1024x8m81_0/wl[82]
+ WL[30] WL[14] bb[14] Cell_array8x8_3v1024x8m81_0/wl[89] WL[31] bb[23] Cell_array8x8_3v1024x8m81_0/wl[92]
+ bb[31] WL[59] Cell_array8x8_3v1024x8m81_0/wl[65] Cell_array8x8_3v1024x8m81_0/wl[75]
+ WL[9] WL[27] WL[34] Cell_array8x8_3v1024x8m81_0/wl[77] Cell_array8x8_3v1024x8m81_0/wl[108]
+ WL[42] Cell_array8x8_3v1024x8m81_0/wl[107] Cell_array8x8_3v1024x8m81_0/wl[78] WL[12]
+ bb[15] Cell_array8x8_3v1024x8m81_0/wl[109] Cell_array8x8_3v1024x8m81_0/wl[112] WL[37]
+ Cell_array8x8_3v1024x8m81_0/wl[111] WL[47] WL[43] Cell_array8x8_3v1024x8m81_0/wl[126]
+ Cell_array8x8_3v1024x8m81_0/wl[81] WL[36] Cell_array8x8_3v1024x8m81_0/wl[98] WL[13]
+ Cell_array8x8_3v1024x8m81_0/wl[100] Cell_array8x8_3v1024x8m81_0/wl[104] WL[22] Cell_array8x8_3v1024x8m81_0/wl[71]
+ Cell_array8x8_3v1024x8m81_0/wl[113] WL[6] bb[7] WL[38] Cell_array8x8_3v1024x8m81_0/wl[99]
+ Cell_array8x8_3v1024x8m81_0/wl[66] WL[20] WL[50] Cell_array8x8_3v1024x8m81_0/wl[114]
+ Cell_array8x8_3v1024x8m81_0/wl[86] Cell_array8x8_3v1024x8m81_0/wl[125] WL[16] Cell_array8x8_3v1024x8m81_0/wl[84]
+ WL[48] Cell_array8x8_3v1024x8m81_0/wl[120] Cell_array8x8_3v1024x8m81_0/wl[83] VDD_uq6
+ WL[35] Cell_array8x8_3v1024x8m81_0/wl[116] WL[33] WL[52] bb[16] Cell_array8x8_3v1024x8m81_0/wl[76]
+ Cell_array8x8_3v1024x8m81_0/wl[85] WL[15] WL[21] WL[49] b[0] WL[127] VSS Cell_array8x8_3v1024x8m81
Xsaout_R_m2_3v1024x8m81_0 ypass[1] ypass[4] ypass[5] saout_m2_3v1024x8m81_4/GWEN din[3]
+ b[0] bb[7] q[3] saout_R_m2_3v1024x8m81_0/vss_uq6 VDD_uq2 VDD_uq0 saout_R_m2_3v1024x8m81_0/vdd_uq2
+ saout_R_m2_3v1024x8m81_0/vdd_uq4 saout_R_m2_3v1024x8m81_0/vdd_uq6 b[1] b[5] bb[6]
+ bb[2] b[7] bb[5] GWE ypass[7] bb[3] WEN[0] bb[0] b[3] saout_R_m2_3v1024x8m81_0/sa_3v1024x8m81_0/pcb
+ men VDD VDD_uq1 b[2] VDD_uq4 VDD_uq3 b[6] bb[4] ypass[3] ypass[2] ypass[6] ypass[0]
+ b[4] VDD_uq5 VSS bb[1] VDD_uq6 saout_R_m2_3v1024x8m81
Xsaout_R_m2_3v1024x8m81_1 ypass[1] ypass[4] ypass[5] saout_m2_3v1024x8m81_4/GWEN din[1]
+ b[16] bb[23] q[1] saout_R_m2_3v1024x8m81_1/vss_uq6 VDD_uq2 VDD_uq0 saout_R_m2_3v1024x8m81_1/vdd_uq2
+ saout_R_m2_3v1024x8m81_1/vdd_uq4 saout_R_m2_3v1024x8m81_1/vdd_uq6 b[17] b[21] bb[22]
+ bb[18] b[23] bb[21] GWE ypass[7] bb[19] WEN[2] bb[16] b[19] saout_R_m2_3v1024x8m81_1/sa_3v1024x8m81_0/pcb
+ men VDD VDD_uq1 b[18] VDD_uq4 VDD_uq3 b[22] bb[20] ypass[3] ypass[2] ypass[6] ypass[0]
+ b[20] VDD_uq5 VSS bb[17] VDD_uq6 saout_R_m2_3v1024x8m81
.ends

.subckt new_dummyrowunit01_3v1024x8m81 018SRAM_cell1_dummy_3v1024x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_2/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_11/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_12/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_3/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_12/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_13/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_4/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_13/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_5/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_14/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_14/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_6/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_15/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_7/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_7/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_8/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_9/m2_134_89# 018SRAM_strap1_3v1024x8m81_1/a_91_178#
+ 018SRAM_cell1_dummy_3v1024x8m81_0/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_0/m2_134_89#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_cell1_dummy_3v1024x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_1/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_10/m2_134_89# VSUBS
X018SRAM_cell1_dummy_3v1024x8m81_10 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_10/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_12 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_12/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_11 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_11/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_13 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_13/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_14 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_14/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_15 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_15/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_0 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_0/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_2 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_2/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_1 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_1/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_3 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_3/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_4 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_4/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_5 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_5/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_6 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_6/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_7 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_7/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_8 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_8/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_9 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_9/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
.ends

.subckt new_dummyrow_unit_3v1024x8m81 018SRAM_cell1_dummy_3v1024x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_2/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_11/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_3/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_12/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_4/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_13/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_14/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_5/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_14/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_6/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_15/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_7/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_7/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_8/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_8/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_9/m2_134_89# 018SRAM_strap1_3v1024x8m81_1/a_91_178#
+ 018SRAM_cell1_dummy_3v1024x8m81_0/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_0/m2_134_89#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_cell1_dummy_3v1024x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_1/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_10/m2_134_89# VSUBS
X018SRAM_cell1_dummy_3v1024x8m81_10 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_10/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_12 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_12/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_11 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_11/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_13 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_13/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_14 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_14/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_15 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_15/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_0 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_0/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_2 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_2/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_1 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_1/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_3 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_3/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_4 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_4/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_5 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_5/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_6 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_6/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_7 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_7/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_8 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_8/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_9 018SRAM_strap1_3v1024x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v1024x8m81_1/w_91_512#
+ 018SRAM_strap1_3v1024x8m81_1/w_91_512# 018SRAM_strap1_3v1024x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v1024x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_9/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
.ends

.subckt x018SRAM_cell1_cutPC_3v1024x8m81 m3_82_330# a_248_342# a_248_592# a_62_178#
+ w_30_512# a_430_96# a_110_96# VSUBS
X0 a_248_592# a_192_298# a_110_250# w_30_512# pfet_03v3 ad=0.1613p pd=1.39u as=0.1238p ps=1.44u w=0.28u l=0.28u
X1 a_248_342# a_192_298# a_110_250# VSUBS nfet_03v3 ad=0.171p pd=1.33u as=0.15665p ps=1.32u w=0.45u l=0.28u
X2 a_192_298# a_110_250# a_248_592# w_30_512# pfet_03v3 ad=0.1238p pd=1.44u as=0.1613p ps=1.39u w=0.28u l=0.28u
X3 a_192_298# a_110_250# a_248_342# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.171p ps=1.33u w=0.45u l=0.28u
X4 a_110_250# a_62_178# a_110_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
X5 a_192_298# a_62_178# a_430_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
.ends

.subckt array16_1024_dummy_01_3v1024x8m81 018SRAM_cell1_cutPC_3v1024x8m81_98/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_81/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_59/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_98/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_59/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_32/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_99/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_106/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_43/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_69/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_91/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_25/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_58/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_69/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_106/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_106/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_98/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_95/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_79/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_102/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_79/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_48/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_21/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_116/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_54/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_87/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_116/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_89/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_89/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_126/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_52/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_109/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_126/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_50/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_5/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_83/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_39/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_99/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_10/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_99/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_10/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_119/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_116/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_1/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_20/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_35/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_68/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_20/a_248_342# VDD_uq0 018SRAM_cell1_cutPC_3v1024x8m81_126/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_107/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_107/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_109/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_30/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_53/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_112/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_37/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_30/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_31/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_64/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_117/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_97/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_117/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_42/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_40/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_40/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_0/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_41/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_127/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_127/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_60/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_93/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_16/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_49/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_32/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_50/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_11/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_50/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_11/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_126/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_5/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_60/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_12/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_21/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_45/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_60/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_78/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_21/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_108/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_108/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_119/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_31/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_70/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_122/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_1/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_52/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_70/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_31/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_71/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_41/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_118/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_74/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_118/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_80/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_41/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_41/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_80/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_115/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_41/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_1/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_61/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_111/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_67/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_107/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_70/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_26/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_59/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_51/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_61/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_73/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_90/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_90/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_12/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_51/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_12/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_121/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_103/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_45/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_83/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_22/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_22/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_61/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_55/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_1/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_61/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_88/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_22/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_109/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_109/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_126/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_71/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_93/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_32/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_51/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_51/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_71/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_32/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_81/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_51/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_84/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_6/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_119/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_119/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_42/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_81/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_2/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_40/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_125/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_81/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_42/a_248_342# VSS_uq0 018SRAM_cell1_cutPC_3v1024x8m81_77/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_117/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_2/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_80/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_36/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_69/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_91/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_13/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_52/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_91/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_52/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_13/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_73/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_113/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_36/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_2/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_62/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_32/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_23/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_65/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_62/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_98/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_23/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_33/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_40/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_72/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_50/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_72/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_33/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_61/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_94/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_17/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_82/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_43/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_39/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_3/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_3/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_82/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_43/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_6/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_127/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_87/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_90/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_13/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_46/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_79/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_92/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_53/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_75/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_92/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_14/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_53/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_14/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_83/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_2/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_123/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_85/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_42/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_63/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_3/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_75/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_24/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_63/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_24/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_100/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_100/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_73/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_95/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_49/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_34/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_73/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_34/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_98/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_108/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_71/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_110/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_27/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_110/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_83/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_4/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_38/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_44/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_4/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_83/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_44/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_120/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_103/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_97/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_104/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_47/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_120/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_23/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_56/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_89/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_93/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_54/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_93/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_15/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_15/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_54/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_113/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_100/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_93/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_50/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_64/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_52/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_4/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_25/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_85/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_7/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_64/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_25/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_123/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_101/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_101/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_74/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_35/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_48/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_74/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_118/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_35/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_81/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_3/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_111/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_37/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_111/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_84/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_37/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_45/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_5/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_67/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_5/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_84/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_45/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_111/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_114/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_121/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_35/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_121/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_33/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_66/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_99/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_94/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_77/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_16/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_55/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_55/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_94/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_16/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_107/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_110/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_39/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_65/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_62/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_5/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_87/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_26/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_95/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_18/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_26/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_65/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_102/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_102/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_103/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_97/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_75/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_36/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_45/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_75/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_7/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_36/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_91/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_112/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_14/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_112/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_47/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_85/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_6/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_36/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_46/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_85/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_6/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_121/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_105/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_122/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_3/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_124/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_122/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_10/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_43/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_76/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_95/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_56/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_95/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_17/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_56/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_17/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_115/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_117/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_120/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_33/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_69/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_109/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_6/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_72/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_66/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_27/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_28/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_66/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_27/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_125/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_103/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_103/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_113/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_76/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_105/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_62/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_47/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_37/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_44/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_37/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_76/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_113/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_24/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_57/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_113/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_7/m3_82_330# VSS VDD 018SRAM_cell1_cutPC_3v1024x8m81_47/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_35/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_69/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_86/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_86/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_7/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_47/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_91/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_123/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_101/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_49/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_123/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_53/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_20/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_86/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_8/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_79/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_96/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_57/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_18/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_57/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_96/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_18/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_127/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_53/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_79/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_119/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_7/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_4/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_82/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_67/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_89/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_38/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_28/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_67/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_28/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_104/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_104/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_123/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_99/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_77/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_75/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_38/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_44/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_115/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_77/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_34/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_38/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_0/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_114/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_34/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_67/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_114/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_8/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_87/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_34/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_48/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_8/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_105/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_87/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_48/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_107/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_124/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_111/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_38/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_124/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_30/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_63/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_96/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_19/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_58/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_97/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_19/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_97/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_58/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_19/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_117/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_42/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_89/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_8/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_92/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_68/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_29/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_15/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_8/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_48/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_68/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_29/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_127/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_105/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_105/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96# 018SRAM_cell1_cutPC_3v1024x8m81_78/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_43/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_85/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_39/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_125/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_4/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_78/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_39/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_11/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_115/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_44/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_77/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_115/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_49/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_88/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_71/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_33/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_88/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_49/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_0/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_121/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_125/m3_82_330# VSUBS 018SRAM_cell1_cutPC_3v1024x8m81_125/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_40/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_73/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_29/a_62_178#
X018SRAM_cell1_cutPC_3v1024x8m81_62 018SRAM_cell1_cutPC_3v1024x8m81_62/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_62/a_248_342# VDD_uq0 018SRAM_cell1_cutPC_3v1024x8m81_62/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_62/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_51 018SRAM_cell1_cutPC_3v1024x8m81_51/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_51/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_51/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_51/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_51/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_40 018SRAM_cell1_cutPC_3v1024x8m81_40/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_40/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_40/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_40/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_40/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_73 018SRAM_cell1_cutPC_3v1024x8m81_73/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_73/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_73/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_73/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_73/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_84 018SRAM_cell1_cutPC_3v1024x8m81_84/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_84/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_87/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_84/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_87/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_95 018SRAM_cell1_cutPC_3v1024x8m81_95/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_95/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_95/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_95/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_95/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_96 018SRAM_cell1_cutPC_3v1024x8m81_96/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_96/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_99/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_96/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_99/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_63 018SRAM_cell1_cutPC_3v1024x8m81_63/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_63/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_2/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_63/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_2/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_52 018SRAM_cell1_cutPC_3v1024x8m81_52/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_52/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_52/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_52/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_52/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_41 018SRAM_cell1_cutPC_3v1024x8m81_41/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_41/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_41/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_41/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_41/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_30 018SRAM_cell1_cutPC_3v1024x8m81_30/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_30/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_32/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_30/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_32/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_74 018SRAM_cell1_cutPC_3v1024x8m81_74/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_74/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_77/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_74/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_77/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_85 018SRAM_cell1_cutPC_3v1024x8m81_85/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_85/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_85/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_85/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_85/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_97 018SRAM_cell1_cutPC_3v1024x8m81_97/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_97/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_97/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_97/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_97/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_31 018SRAM_cell1_cutPC_3v1024x8m81_31/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_31/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_61/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_31/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_61/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_53 018SRAM_cell1_cutPC_3v1024x8m81_53/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_53/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_53/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_53/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_53/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_20 018SRAM_cell1_cutPC_3v1024x8m81_20/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_20/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_42/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_20/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_42/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_42 018SRAM_cell1_cutPC_3v1024x8m81_42/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_42/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_42/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_42/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_42/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_64 018SRAM_cell1_cutPC_3v1024x8m81_64/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_64/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_67/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_64/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_67/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_75 018SRAM_cell1_cutPC_3v1024x8m81_75/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_75/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_75/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_75/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_75/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_86 018SRAM_cell1_cutPC_3v1024x8m81_86/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_86/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_89/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_86/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_89/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_98 018SRAM_cell1_cutPC_3v1024x8m81_98/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_98/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_98/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_98/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_98/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_54 018SRAM_cell1_cutPC_3v1024x8m81_54/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_54/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_54/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_9/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_10 018SRAM_cell1_cutPC_3v1024x8m81_10/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_10/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_53/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_10/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_53/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_43 018SRAM_cell1_cutPC_3v1024x8m81_43/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_43/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_43/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_43/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_43/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_21 018SRAM_cell1_cutPC_3v1024x8m81_21/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_21/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_41/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_21/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_41/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_32 018SRAM_cell1_cutPC_3v1024x8m81_32/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_32/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_32/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_32/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_32/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_65 018SRAM_cell1_cutPC_3v1024x8m81_65/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_65/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_1/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_65/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_76 018SRAM_cell1_cutPC_3v1024x8m81_76/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_76/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_79/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_76/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_79/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_87 018SRAM_cell1_cutPC_3v1024x8m81_87/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_87/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_87/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_87/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_87/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_99 018SRAM_cell1_cutPC_3v1024x8m81_99/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_99/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_99/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_99/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_99/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_55 018SRAM_cell1_cutPC_3v1024x8m81_55/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_55/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_8/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_55/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_8/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_11 018SRAM_cell1_cutPC_3v1024x8m81_11/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_11/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_52/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_11/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_52/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_44 018SRAM_cell1_cutPC_3v1024x8m81_44/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_44/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_44/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_44/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_44/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_22 018SRAM_cell1_cutPC_3v1024x8m81_22/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_22/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_40/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_22/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_40/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_33 018SRAM_cell1_cutPC_3v1024x8m81_33/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_33/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_33/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_33/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_33/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_66 018SRAM_cell1_cutPC_3v1024x8m81_66/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_66/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_69/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_66/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_69/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_77 018SRAM_cell1_cutPC_3v1024x8m81_77/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_77/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_77/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_77/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_77/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_88 018SRAM_cell1_cutPC_3v1024x8m81_88/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_88/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_91/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_88/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_91/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_56 018SRAM_cell1_cutPC_3v1024x8m81_56/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_56/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_7/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_56/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_7/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_12 018SRAM_cell1_cutPC_3v1024x8m81_12/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_12/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_51/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_12/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_51/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_45 018SRAM_cell1_cutPC_3v1024x8m81_45/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_45/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_45/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_45/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_45/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_23 018SRAM_cell1_cutPC_3v1024x8m81_23/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_23/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_39/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_23/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_39/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_34 018SRAM_cell1_cutPC_3v1024x8m81_34/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_34/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_34/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_34/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_34/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_67 018SRAM_cell1_cutPC_3v1024x8m81_67/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_67/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_67/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_67/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_67/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_78 018SRAM_cell1_cutPC_3v1024x8m81_78/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_78/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_81/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_78/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_81/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_89 018SRAM_cell1_cutPC_3v1024x8m81_89/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_89/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_89/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_89/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_89/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_57 018SRAM_cell1_cutPC_3v1024x8m81_57/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_57/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_6/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_57/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_6/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_13 018SRAM_cell1_cutPC_3v1024x8m81_13/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_13/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_50/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_13/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_50/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_46 018SRAM_cell1_cutPC_3v1024x8m81_46/m3_82_330#
+ VSS VDD 018SRAM_cell1_cutPC_3v1024x8m81_46/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_24 018SRAM_cell1_cutPC_3v1024x8m81_24/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_24/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_38/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_24/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_38/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_35 018SRAM_cell1_cutPC_3v1024x8m81_35/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_35/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_35/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_35/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_35/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_68 018SRAM_cell1_cutPC_3v1024x8m81_68/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_68/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_71/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_68/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_71/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_79 018SRAM_cell1_cutPC_3v1024x8m81_79/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_79/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_79/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_79/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_79/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_58 018SRAM_cell1_cutPC_3v1024x8m81_58/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_58/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_5/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_58/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_5/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_14 018SRAM_cell1_cutPC_3v1024x8m81_14/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_14/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_49/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_14/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_49/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_0 018SRAM_cell1_cutPC_3v1024x8m81_0/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_0/a_248_342#
+ VDD 018SRAM_cell1_cutPC_3v1024x8m81_0/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_0/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_47 018SRAM_cell1_cutPC_3v1024x8m81_47/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_47/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_47/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_47/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_47/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_25 018SRAM_cell1_cutPC_3v1024x8m81_25/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_25/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_37/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_25/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_37/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_36 018SRAM_cell1_cutPC_3v1024x8m81_36/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_36/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_36/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_36/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_36/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_69 018SRAM_cell1_cutPC_3v1024x8m81_69/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_69/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_69/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_69/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_69/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_59 018SRAM_cell1_cutPC_3v1024x8m81_59/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_59/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_4/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_59/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_4/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_15 018SRAM_cell1_cutPC_3v1024x8m81_15/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_15/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_48/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_15/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_48/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_48 018SRAM_cell1_cutPC_3v1024x8m81_48/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_48/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_48/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_48/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_48/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_37 018SRAM_cell1_cutPC_3v1024x8m81_37/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_37/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_37/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_37/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_37/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_26 018SRAM_cell1_cutPC_3v1024x8m81_26/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_26/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_36/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_26/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_36/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_1 018SRAM_cell1_cutPC_3v1024x8m81_1/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_1/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_1/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_1/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_120 018SRAM_cell1_cutPC_3v1024x8m81_120/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_120/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_123/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_120/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_123/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_2 018SRAM_cell1_cutPC_3v1024x8m81_2/m3_82_330# VSS_uq0
+ 018SRAM_cell1_cutPC_3v1024x8m81_2/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_2/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_2/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_16 018SRAM_cell1_cutPC_3v1024x8m81_16/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_16/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_45/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_16/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_45/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_121 018SRAM_cell1_cutPC_3v1024x8m81_121/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_121/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_121/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_121/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_121/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_110 018SRAM_cell1_cutPC_3v1024x8m81_110/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_110/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_113/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_110/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_113/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_49 018SRAM_cell1_cutPC_3v1024x8m81_49/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_49/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_49/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_49/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_49/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_38 018SRAM_cell1_cutPC_3v1024x8m81_38/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_38/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_38/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_38/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_38/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_27 018SRAM_cell1_cutPC_3v1024x8m81_27/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_27/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_35/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_27/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_35/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_3 018SRAM_cell1_cutPC_3v1024x8m81_3/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_3/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_3/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_3/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_3/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_17 018SRAM_cell1_cutPC_3v1024x8m81_17/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_17/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_47/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_17/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_47/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_39 018SRAM_cell1_cutPC_3v1024x8m81_39/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_39/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_39/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_39/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_39/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_28 018SRAM_cell1_cutPC_3v1024x8m81_28/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_28/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_34/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_28/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_34/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_122 018SRAM_cell1_cutPC_3v1024x8m81_122/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_122/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_125/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_122/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_125/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_111 018SRAM_cell1_cutPC_3v1024x8m81_111/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_111/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_111/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_111/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_111/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_100 018SRAM_cell1_cutPC_3v1024x8m81_100/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_100/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_103/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_100/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_103/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_4 018SRAM_cell1_cutPC_3v1024x8m81_4/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_4/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_4/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_4/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_4/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_123 018SRAM_cell1_cutPC_3v1024x8m81_123/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_123/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_123/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_123/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_123/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_112 018SRAM_cell1_cutPC_3v1024x8m81_112/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_112/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_115/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_112/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_115/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_101 018SRAM_cell1_cutPC_3v1024x8m81_101/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_101/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_98/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_101/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_98/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_18 018SRAM_cell1_cutPC_3v1024x8m81_18/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_18/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_44/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_18/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_44/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_29 018SRAM_cell1_cutPC_3v1024x8m81_29/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_29/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_33/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_29/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_33/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_5 018SRAM_cell1_cutPC_3v1024x8m81_5/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_5/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_5/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_5/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_5/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_19 018SRAM_cell1_cutPC_3v1024x8m81_19/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_19/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_43/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_19/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_43/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_124 018SRAM_cell1_cutPC_3v1024x8m81_124/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_124/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_127/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_124/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_127/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_113 018SRAM_cell1_cutPC_3v1024x8m81_113/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_113/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_113/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_113/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_113/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_102 018SRAM_cell1_cutPC_3v1024x8m81_102/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_102/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_105/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_102/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_105/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_6 018SRAM_cell1_cutPC_3v1024x8m81_6/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_6/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_6/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_6/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_6/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_125 018SRAM_cell1_cutPC_3v1024x8m81_125/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_125/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_125/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_125/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_125/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_114 018SRAM_cell1_cutPC_3v1024x8m81_114/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_114/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_117/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_114/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_117/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_103 018SRAM_cell1_cutPC_3v1024x8m81_103/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_103/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_103/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_103/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_103/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_7 018SRAM_cell1_cutPC_3v1024x8m81_7/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_7/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_7/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_7/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_7/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_126 018SRAM_cell1_cutPC_3v1024x8m81_126/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_126/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_126/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_126/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_126/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_115 018SRAM_cell1_cutPC_3v1024x8m81_115/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_115/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_115/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_115/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_115/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_104 018SRAM_cell1_cutPC_3v1024x8m81_104/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_104/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_107/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_104/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_107/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_8 018SRAM_cell1_cutPC_3v1024x8m81_8/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_8/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_8/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_8/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_8/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_116 018SRAM_cell1_cutPC_3v1024x8m81_116/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_116/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_119/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_116/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_119/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_105 018SRAM_cell1_cutPC_3v1024x8m81_105/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_105/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_105/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_105/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_105/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_127 018SRAM_cell1_cutPC_3v1024x8m81_127/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_127/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_127/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_127/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_127/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_9 018SRAM_cell1_cutPC_3v1024x8m81_9/m3_82_330# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_248_342#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_248_592# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_62_178#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/w_30_512# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_117 018SRAM_cell1_cutPC_3v1024x8m81_117/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_117/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_117/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_117/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_117/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_106 018SRAM_cell1_cutPC_3v1024x8m81_106/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_106/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_109/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_106/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_109/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_118 018SRAM_cell1_cutPC_3v1024x8m81_118/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_118/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_121/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_118/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_121/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_107 018SRAM_cell1_cutPC_3v1024x8m81_107/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_107/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_107/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_107/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_107/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_119 018SRAM_cell1_cutPC_3v1024x8m81_119/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_119/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_119/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_119/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_119/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_108 018SRAM_cell1_cutPC_3v1024x8m81_108/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_108/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_111/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_108/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_111/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_109 018SRAM_cell1_cutPC_3v1024x8m81_109/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_109/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_109/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_109/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_109/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_90 018SRAM_cell1_cutPC_3v1024x8m81_90/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_90/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_93/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_90/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_93/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_80 018SRAM_cell1_cutPC_3v1024x8m81_80/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_80/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_83/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_80/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_83/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_91 018SRAM_cell1_cutPC_3v1024x8m81_91/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_91/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_91/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_91/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_91/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_70 018SRAM_cell1_cutPC_3v1024x8m81_70/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_70/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_73/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_70/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_73/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_81 018SRAM_cell1_cutPC_3v1024x8m81_81/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_81/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_81/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_81/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_81/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_92 018SRAM_cell1_cutPC_3v1024x8m81_92/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_92/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_95/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_92/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_95/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_60 018SRAM_cell1_cutPC_3v1024x8m81_60/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_60/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_3/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_60/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_3/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_71 018SRAM_cell1_cutPC_3v1024x8m81_71/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_71/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_71/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_71/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_71/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_82 018SRAM_cell1_cutPC_3v1024x8m81_82/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_82/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_85/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_82/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_85/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_93 018SRAM_cell1_cutPC_3v1024x8m81_93/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_93/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_93/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_93/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_93/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_61 018SRAM_cell1_cutPC_3v1024x8m81_61/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_61/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_61/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_61/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_61/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_50 018SRAM_cell1_cutPC_3v1024x8m81_50/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_50/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_50/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_50/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_50/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_72 018SRAM_cell1_cutPC_3v1024x8m81_72/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_72/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_75/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_72/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_75/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_83 018SRAM_cell1_cutPC_3v1024x8m81_83/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_83/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_83/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_83/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_83/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
X018SRAM_cell1_cutPC_3v1024x8m81_94 018SRAM_cell1_cutPC_3v1024x8m81_94/m3_82_330#
+ 018SRAM_cell1_cutPC_3v1024x8m81_94/a_248_342# 018SRAM_cell1_cutPC_3v1024x8m81_97/a_248_592#
+ 018SRAM_cell1_cutPC_3v1024x8m81_94/a_62_178# 018SRAM_cell1_cutPC_3v1024x8m81_97/w_30_512#
+ 018SRAM_cell1_cutPC_3v1024x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v1024x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v1024x8m81
.ends

.subckt ldummy_3v512x4_3v1024x8m81 018SRAM_cell1_dummy_3v1024x8m81_30/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_83/a_248_592#
+ 018SRAM_cell1_dummy_3v1024x8m81_30/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_61/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_22/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_61/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_22/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_10/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_116/m3_82_330#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_10/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_116/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_42/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_89/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_71/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_93/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_8/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_32/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_51/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_71/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_32/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_126/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_109/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_126/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_2/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_11/m2_346_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_85/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_81/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_2/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_11/m2_134_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_42/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_40/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_125/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_42/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_81/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_119/a_248_592#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_5/m2_346_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_5/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_21/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_9/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_91/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_52/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_21/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_13/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_9/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_91/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_52/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_13/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_107/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_107/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_31/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_62/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_23/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_31/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_62/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_6/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_23/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_11/m2_346_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_10/m2_346_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_117/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_117/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_11/m2_134_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_10/m2_134_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_32/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_99/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_43/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_9/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_72/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_50/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_33/m3_82_330#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_0/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_72/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_33/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_127/m3_82_330#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_0/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_2/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_127/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_3/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_12/m2_346_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_82/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_3/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_12/m2_134_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_43/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_95/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_39/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_82/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_48/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_43/a_248_342#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_6/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_22/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_6/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_92/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_75/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_14/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_53/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_22/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_92/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_53/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_14/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_52/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_108/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_108/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_63/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_85/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_24/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_63/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_24/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_12/m2_346_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_11/m2_346_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_118/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_118/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_12/m2_134_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_11/m2_134_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_95/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_49/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_73/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_34/m3_82_330#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_1/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_73/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_34/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_111/a_248_592#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_1/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_4/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_83/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_4/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_37/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_38/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_44/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_13/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_83/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_44/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_121/a_248_592#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_7/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/VSS
+ array16_1024_dummy_01_3v1024x8m81_0/VDD new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_7/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_23/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_0/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_93/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_54/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_23/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_93/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_15/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_0/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_54/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_41/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_15/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_109/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_109/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_25/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_64/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_64/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_13/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_25/a_248_342#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_12/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_119/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_119/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_13/m2_134_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_12/m2_134_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_74/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_35/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_48/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_74/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_2/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_35/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_2/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_14/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_5/m2_134_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_37/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_45/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_14/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_84/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_67/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_84/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_71/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_45/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_111/w_30_512#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_8/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_24/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_8/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_7/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_94/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_77/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_1/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_16/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_55/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_24/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_55/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_94/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_16/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_61/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_67/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_107/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_65/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_87/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_26/m3_82_330#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_14/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_3/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_65/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_26/a_248_342#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_13/m2_346_89# new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_14/m2_134_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_13/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_103/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_45/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_97/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_1/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_75/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_36/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_75/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_45/a_248_592#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_3/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_36/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_3/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_15/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_85/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_6/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_51/w_30_512#
+ 018SRAM_cell1_dummy_3v1024x8m81_15/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_36/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_46/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_85/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_81/w_30_512#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_9/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_25/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_9/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_2/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_56/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_95/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_25/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_95/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_17/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_56/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_17/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_100/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_77/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_117/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_100/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_66/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_27/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_66/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_15/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_27/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_110/m3_82_330#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_14/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_110/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_15/m2_134_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_14/m2_134_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_73/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_113/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_36/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_2/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_76/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_47/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_37/m3_82_330#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_4/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_76/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_37/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_120/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_103/a_248_592#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_4/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_120/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_7/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_16/m2_346_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_40/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_47/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_69/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_86/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_7/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_16/m2_134_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_35/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_86/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_47/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_113/a_248_592#
+ 018SRAM_cell1_dummy_3v1024x8m81_26/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_3/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_79/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_96/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_3/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_26/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_57/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_18/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_96/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_57/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_18/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_123/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_101/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_87/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_101/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_127/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_67/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_89/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_28/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_67/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_28/a_248_342#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_15/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_111/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_111/a_248_342#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_15/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_83/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_123/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_3/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_99/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_77/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_38/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_44/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_38/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_5/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_77/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_121/m3_82_330#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_5/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_121/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_8/w_30_512#
+ 018SRAM_cell1_dummy_3v1024x8m81_8/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_17/m2_346_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_87/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_8/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_34/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_48/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_17/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_98/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_87/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_48/a_248_342#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_0/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_27/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_0/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_4/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_4/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_58/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_97/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_4/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_27/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_19/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_97/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_58/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_19/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_97/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_102/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_47/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_102/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_68/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_0/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_29/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_29/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_68/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_112/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_112/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_93/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_50/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_4/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_78/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_43/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_39/m3_82_330#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_6/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_78/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_39/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_105/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_122/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_122/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_6/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_18/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_9/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_9/m2_134_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_88/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_71/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_33/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_49/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_18/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_88/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_49/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_115/a_248_592#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_1/m2_346_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_1/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_28/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_98/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_5/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_59/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_28/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_81/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_5/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_98/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_59/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_125/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_103/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_103/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_35/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_69/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_91/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_69/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_113/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_113/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_39/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_5/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_98/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_79/m3_82_330#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_7/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_79/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_123/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_123/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_7/m2_134_89# 018SRAM_cell1_dummy_3v1024x8m81_19/m2_346_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_89/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_19/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_89/a_248_342#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_2/m2_346_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_2/m2_134_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_29/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_6/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_99/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_6/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_10/m3_82_330#
+ 018SRAM_cell1_dummy_3v1024x8m81_29/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_99/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_10/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_104/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_121/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_104/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_20/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_20/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_9/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_114/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_114/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_33/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_69/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_109/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_6/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_30/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_53/a_248_592#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_8/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_30/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_107/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_124/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_124/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_8/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_5/w_30_512#
+ 018SRAM_cell1_dummy_3v1024x8m81_0/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_0/m2_134_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_40/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_105/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_42/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_44/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_40/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_117/a_248_592#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_3/m2_346_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_3/m2_134_89#
+ array16_1024_dummy_01_3v1024x8m81_0/VSS_uq0 array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_1/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_7/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_32/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_50/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_11/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_7/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_50/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_11/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_91/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_127/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_49/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_105/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_105/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_60/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_21/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_60/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_21/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_115/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_115/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_53/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_79/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_119/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_7/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_31/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_70/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_52/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_31/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_70/a_248_342#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_9/m2_346_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_125/m3_82_330#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_9/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_125/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_1/m2_346_89# 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_3v1024x8m81_10/m2_346_89# m3_5692_40200# 018SRAM_cell1_dummy_3v1024x8m81_1/m2_134_89#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_80/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_75/w_30_512#
+ 018SRAM_cell1_dummy_3v1024x8m81_10/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_41/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_41/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_34/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_80/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_115/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_41/a_248_342#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_4/m2_346_89# 018SRAM_cell1_dummy_3v1024x8m81_20/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_4/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_8/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_51/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_73/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_90/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_8/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_90/a_248_342#
+ 018SRAM_cell1_dummy_3v1024x8m81_20/m2_134_89# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_61/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_12/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_51/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_12/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_38/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_106/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_106/a_248_342#
X018SRAM_cell1_3v1024x8m81_1 VSUBS VSUBS 018SRAM_cell1_3v1024x8m81_1/w_30_512# VSUBS
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# 018SRAM_cell1_3v1024x8m81_1/a_430_96# 018SRAM_cell1_3v1024x8m81_1/a_110_96#
+ VSUBS x018SRAM_cell1_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_30 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_30/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_30/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_20 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_20/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_20/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_31 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_31/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_31/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_21 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_21/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_21/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_10 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_10/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_22 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_22/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_22/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_11 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_11/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_23 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_23/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_23/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_12 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_12/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_24 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_24/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_24/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_13 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_13/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
Xnew_dummyrowunit01_3v1024x8m81_0 new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_2/m2_346_89#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_2/m2_134_89# new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_11/m2_346_89#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_11/m2_134_89# new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_3/m2_346_89#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_12/m2_134_89# new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_3/m2_134_89#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_12/m2_346_89# new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_4/m2_346_89#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_13/m2_134_89# new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_4/m2_134_89#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_13/m2_346_89# new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_5/m2_346_89#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_5/m2_134_89# new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_14/m2_134_89#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_14/m2_346_89# new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_6/m2_346_89#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_6/m2_134_89# new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_15/m2_346_89#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_15/m2_134_89# new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_7/m2_134_89#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_7/m2_346_89# new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_8/m2_346_89#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_8/m2_134_89# new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_9/m2_346_89#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_9/m2_134_89# VSUBS
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_0/m2_346_89# new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_0/m2_134_89#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_1/m2_346_89#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_1/m2_134_89# new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_10/m2_346_89#
+ new_dummyrowunit01_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_10/m2_134_89# VSUBS
+ new_dummyrowunit01_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_25 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_25/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_25/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_14 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_14/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_15 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_15/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_26 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_26/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_26/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_27 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_27/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_27/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_16 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_16/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_16/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_28 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_28/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_28/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_17 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_17/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_17/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_29 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_29/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_29/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_18 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_18/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_18/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_19 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_19/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_19/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_0 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_0/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
Xnew_dummyrow_unit_3v1024x8m81_0 new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_2/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_2/m2_134_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_11/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_11/m2_134_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_3/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_3/m2_134_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_12/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_12/m2_134_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_4/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_4/m2_134_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_13/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_13/m2_134_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_5/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_14/m2_134_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_5/m2_134_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_14/m2_346_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_6/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_6/m2_134_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_15/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_15/m2_134_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_7/m2_134_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_7/m2_346_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_8/m2_134_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_8/m2_346_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_9/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_9/m2_134_89# VSUBS
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_0/m2_346_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_0/m2_134_89#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_1/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_1/m2_134_89# new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_10/m2_346_89#
+ new_dummyrow_unit_3v1024x8m81_0/018SRAM_cell1_dummy_3v1024x8m81_10/m2_134_89# VSUBS
+ new_dummyrow_unit_3v1024x8m81
Xarray16_1024_dummy_01_3v1024x8m81_0 array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_98/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_81/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_59/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_98/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_59/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_32/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_99/w_30_512#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_43/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_9/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_69/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_91/a_248_592#
+ VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_69/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_106/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_106/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_98/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_95/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_79/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_79/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_48/w_30_512#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_116/m3_82_330#
+ VSUBS VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_116/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_89/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_89/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_126/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_52/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_109/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_126/a_248_342#
+ VSUBS VSUBS VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_99/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_10/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_99/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_10/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_119/a_248_592#
+ VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_20/m3_82_330#
+ VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_20/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 018SRAM_cell1_3v1024x8m81_1/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_107/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_107/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_109/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_30/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_53/a_248_592#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_37/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_30/a_248_342#
+ VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_117/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_117/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_42/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_0/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_40/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_40/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_0/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_41/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_127/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_9/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_127/a_248_342#
+ VSUBS VSUBS VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_32/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_50/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_11/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_50/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_11/a_248_342#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_5/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_60/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_21/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_60/a_248_342#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_21/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_108/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_108/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_119/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_31/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_70/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_1/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_52/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_70/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_31/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_71/w_30_512#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_118/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_118/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_80/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_1/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_41/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_41/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_80/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_115/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_41/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_1/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_61/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_111/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_67/w_30_512#
+ VSUBS VSUBS VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_51/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_61/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_73/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_90/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_90/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_12/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_51/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_12/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_121/a_248_592#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_45/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_83/a_248_592#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_22/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_61/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_1/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_61/a_248_342#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_22/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_109/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_109/a_248_342#
+ 018SRAM_cell1_3v1024x8m81_1/w_30_512# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_71/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_93/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_32/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_51/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_51/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_71/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_32/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_81/w_30_512#
+ VSUBS VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_119/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_119/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_42/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_81/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_2/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_40/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_125/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_81/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_42/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/VSS_uq0 array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_77/w_30_512#
+ VSUBS VSUBS VSUBS VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_91/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_13/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_52/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_91/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_52/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_13/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_73/w_30_512#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_36/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_2/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_62/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_23/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_62/a_248_342#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_23/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_33/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_40/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_72/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_50/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_72/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_33/a_248_342#
+ VSUBS VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_82/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_43/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_39/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_3/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_3/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_82/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_43/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_6/w_30_512#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_87/w_30_512#
+ VSUBS VSUBS VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_92/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_53/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_75/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_92/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_14/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_53/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_14/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_83/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_2/w_30_512#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_85/a_248_592#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_63/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_3/a_248_592#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_24/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_63/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_24/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_100/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_100/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_73/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_95/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_49/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_34/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_73/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_34/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_98/w_30_512#
+ VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_110/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_110/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_83/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_4/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_38/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_44/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_4/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_83/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_44/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_120/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_103/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_97/w_30_512#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_47/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_120/a_248_342#
+ VSUBS VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_93/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_54/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_93/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_15/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_15/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_54/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_113/a_248_592#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_93/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_50/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_64/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_4/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_25/m3_82_330#
+ VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_64/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_25/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_123/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_101/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_101/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_74/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_35/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_48/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_74/a_248_342#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_35/a_248_342#
+ VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_111/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_111/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_84/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_37/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_45/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_5/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_67/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_5/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_84/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_45/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_111/w_30_512#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_121/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_35/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_121/a_248_342#
+ VSUBS VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_94/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_77/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_16/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_55/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_55/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_94/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_16/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_107/w_30_512#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_39/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_65/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_5/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_87/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_26/m3_82_330#
+ VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_26/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_65/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_102/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_102/a_248_342#
+ 018SRAM_cell1_3v1024x8m81_1/a_430_96# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_103/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_97/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_75/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_36/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_45/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_75/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_7/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_36/a_248_342#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_112/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_112/a_248_342#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_85/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_6/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_36/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_46/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_85/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_6/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_121/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_105/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_122/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_3/w_30_512#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_122/a_248_342#
+ VSUBS VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_95/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_56/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_95/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_17/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_56/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_17/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_115/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_117/w_30_512#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_33/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_69/w_30_512#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_6/a_248_592#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_66/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_27/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_66/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_27/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_125/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_103/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_103/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_113/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_76/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_47/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_37/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_44/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_37/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_76/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_113/m3_82_330#
+ VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_113/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_7/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/VSS array16_1024_dummy_01_3v1024x8m81_0/VDD
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_47/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_35/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_69/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_86/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_86/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_7/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_47/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_91/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_123/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_49/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_123/a_248_342#
+ VSUBS VSUBS VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_79/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_96/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_57/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_18/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_57/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_96/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_18/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_127/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_53/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_79/w_30_512#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_7/a_248_592#
+ VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_67/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_89/a_248_592#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_28/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_67/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_28/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_104/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_104/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_123/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_99/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_77/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_75/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_38/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_44/a_248_592#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_77/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_34/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_38/a_248_342#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_114/m3_82_330#
+ VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_114/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_8/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_87/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_34/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_48/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_8/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_105/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_87/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_48/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_107/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_124/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_38/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_124/a_248_342#
+ VSUBS VSUBS VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_58/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_97/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_19/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_97/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_58/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_19/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_117/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_42/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_89/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_8/w_30_512#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_68/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_29/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_8/a_248_592#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_68/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_29/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_127/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_105/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_105/a_248_342#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_78/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_43/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_85/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_39/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_4/w_30_512#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_78/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_39/a_248_342#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_115/m3_82_330#
+ VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_115/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_9/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_49/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_88/m3_82_330#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_71/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_33/a_248_592#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_88/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_9/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_49/a_248_342#
+ array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_0/w_30_512#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_125/m3_82_330#
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/018SRAM_cell1_cutPC_3v1024x8m81_125/a_248_342#
+ VSUBS VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_1 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_1/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_2 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_2/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_3 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_3/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_4 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_4/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_5 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_5/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_6 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_6/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_7 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_7/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_8 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_8/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_dummy_3v1024x8m81_9 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v1024x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v1024x8m81_9/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v1024x8m81
X018SRAM_cell1_3v1024x8m81_0 VSUBS VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0
+ VSUBS array16_1024_dummy_01_3v1024x8m81_0/VDD_uq0 018SRAM_cell1_3v1024x8m81_1/a_430_96#
+ 018SRAM_cell1_3v1024x8m81_1/a_110_96# VSUBS x018SRAM_cell1_3v1024x8m81
.ends

.subckt lcol4_1024_3v1024x8m81 WL[32] WL[33] WL[34] WL[38] WL[39] WL[35] WL[36] WL[37]
+ WL[41] WL[43] WL[45] WL[48] WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56]
+ WL[58] WL[60] WL[63] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12]
+ WL[10] WL[9] WL[8] WL[6] WL[31] WL[30] WL[29] din[1] din[3] din[2] q[1] q[2] q[3]
+ pcb[2] pcb[3] pcb[0] pcb[1] WEN[3] WEN[2] WEN[1] q[0] d[0] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[76]
+ col_1024a_3v1024x8m81_0/WL[14] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[113]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[86] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[123]
+ col_1024a_3v1024x8m81_0/WL[15] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[96]
+ col_1024a_3v1024x8m81_0/WL[32] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[69]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[102] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[79]
+ col_1024a_3v1024x8m81_0/WL[17] col_1024a_3v1024x8m81_0/WL[34] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[112]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[89] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[122]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[99] col_1024a_3v1024x8m81_0/WL[19]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[68] col_1024a_3v1024x8m81_0/WL[36]
+ col_1024a_3v1024x8m81_0/saout_R_m2_3v1024x8m81_0/vdd_uq4 col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[105]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[78] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[115]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[88] col_1024a_3v1024x8m81_0/WL[38]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[125] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[98]
+ col_1024a_3v1024x8m81_0/WL[39] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[104]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[114] col_1024a_3v1024x8m81_0/WL[58]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[124] WL[57] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[107]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[71] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[117]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[81] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[91]
+ col_1024a_3v1024x8m81_0/saout_m2_3v1024x8m81_4/GWEN col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[106]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[70] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[116]
+ col_1024a_3v1024x8m81_0/WL[21] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[80]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[126] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[90]
+ WL[21] col_1024a_3v1024x8m81_0/ypass[0] WL[22] col_1024a_3v1024x8m81_0/WL[40] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[109]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[73] col_1024a_3v1024x8m81_0/ypass[1]
+ WL[23] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[119] col_1024a_3v1024x8m81_0/WL[41]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[83] col_1024a_3v1024x8m81_0/ypass[2]
+ WL[24] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[93] WL[40] col_1024a_3v1024x8m81_0/ypass[3]
+ WL[25] col_1024a_3v1024x8m81_0/WL[43] col_1024a_3v1024x8m81_0/WL[60] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[108]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[72] col_1024a_3v1024x8m81_0/ypass[4]
+ WL[26] WL[42] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[118] WL[59]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[82] col_1024a_3v1024x8m81_0/ypass[5]
+ WL[27] col_1024a_3v1024x8m81_0/WL[45] col_1024a_3v1024x8m81_0/WL[62] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[92]
+ col_1024a_3v1024x8m81_0/ypass[6] WL[28] WL[44] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[65]
+ col_1024a_3v1024x8m81_0/ypass[7] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[75]
+ col_1024a_3v1024x8m81_0/WL[47] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[85]
+ col_1024a_3v1024x8m81_0/VDD_uq5 col_1024a_3v1024x8m81_0/WL[127] WL[46] WL[0] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[95]
+ col_1024a_3v1024x8m81_0/VDD_uq4 WL[47] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[64]
+ WL[1] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[101] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[74]
+ WL[2] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[111] col_1024a_3v1024x8m81_0/VDD_uq2
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[84] WL[3] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[121]
+ col_1024a_3v1024x8m81_0/VDD_uq1 col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[94]
+ WL[4] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[67] WL[61] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[100]
+ col_1024a_3v1024x8m81_0/WL[10] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[77]
+ WL[5] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[110] WL[11] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[87]
+ col_1024a_3v1024x8m81_0/VDD_uq3 col_1024a_3v1024x8m81_0/WL[6] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[120]
+ WEN[0] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[97] col_1024a_3v1024x8m81_0/WL[12]
+ WL[7] col_1024a_3v1024x8m81_0/VDD_uq0 col_1024a_3v1024x8m81_0/GWE col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[66]
+ col_1024a_3v1024x8m81_0/men VDD col_1024a_3v1024x8m81_0/WL[13] col_1024a_3v1024x8m81_0/VDD
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[103] col_1024a_3v1024x8m81_0/WL[8]
+ VSUBS
Xcol_1024a_3v1024x8m81_0 WL[3] col_1024a_3v1024x8m81_0/ypass[0] col_1024a_3v1024x8m81_0/ypass[1]
+ col_1024a_3v1024x8m81_0/ypass[3] col_1024a_3v1024x8m81_0/ypass[4] col_1024a_3v1024x8m81_0/ypass[5]
+ col_1024a_3v1024x8m81_0/VDD col_1024a_3v1024x8m81_0/WL[32] WL[30] WL[29] WL[22]
+ WL[21] WL[55] WL[19] WL[46] col_1024a_3v1024x8m81_0/WL[12] WL[11] WL[48] WL[49]
+ col_1024a_3v1024x8m81_0/WL[41] col_1024a_3v1024x8m81_0/WL[40] col_1024a_3v1024x8m81_0/WL[10]
+ col_1024a_3v1024x8m81_0/WL[43] WL[34] col_1024a_3v1024x8m81_0/WL[34] WL[36] WL[32]
+ col_1024a_3v1024x8m81_0/WL[38] col_1024a_3v1024x8m81_0/WL[36] WL[5] WL[17] WL[53]
+ WL[51] col_1024a_3v1024x8m81_0/WL[17] WL[52] WL[50] col_1024a_3v1024x8m81_0/WL[127]
+ WL[59] col_1024a_3v1024x8m81_0/WL[15] col_1024a_3v1024x8m81_0/WL[14] col_1024a_3v1024x8m81_0/WL[13]
+ WL[0] col_1024a_3v1024x8m81_0/ypass[2] WL[24] col_1024a_3v1024x8m81_0/b[16] col_1024a_3v1024x8m81_0/b[19]
+ din[1] din[3] din[2] d[0] q[0] q[1] q[2] q[3] col_1024a_3v1024x8m81_0/b[17] col_1024a_3v1024x8m81_0/b[14]
+ col_1024a_3v1024x8m81_0/b[8] col_1024a_3v1024x8m81_0/bb[8] col_1024a_3v1024x8m81_0/bb[10]
+ col_1024a_3v1024x8m81_0/bb[11] col_1024a_3v1024x8m81_0/bb[12] col_1024a_3v1024x8m81_0/bb[13]
+ col_1024a_3v1024x8m81_0/bb[14] col_1024a_3v1024x8m81_0/bb[15] col_1024a_3v1024x8m81_0/bb[16]
+ col_1024a_3v1024x8m81_0/bb[24] col_1024a_3v1024x8m81_0/bb[25] col_1024a_3v1024x8m81_0/bb[27]
+ col_1024a_3v1024x8m81_0/bb[29] col_1024a_3v1024x8m81_0/bb[30] col_1024a_3v1024x8m81_0/bb[31]
+ col_1024a_3v1024x8m81_0/b[30] col_1024a_3v1024x8m81_0/b[24] col_1024a_3v1024x8m81_0/b[0]
+ col_1024a_3v1024x8m81_0/b[18] col_1024a_3v1024x8m81_0/pcb[0] col_1024a_3v1024x8m81_0/pcb[1]
+ col_1024a_3v1024x8m81_0/pcb[3] col_1024a_3v1024x8m81_0/pcb[2] WEN[3] WEN[2] WEN[0]
+ col_1024a_3v1024x8m81_0/VDD_uq5 col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[81]
+ col_1024a_3v1024x8m81_0/WL[39] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[108]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[126] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[75]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[93] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[111]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[70] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/b[8]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[88] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[90]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[124] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[73]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[91] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[118]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[109] col_1024a_3v1024x8m81_0/ypass[6]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[68] col_1024a_3v1024x8m81_0/ypass[7]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[86] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[104]
+ VSUBS col_1024a_3v1024x8m81_0/men col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[71]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[98] WL[1] col_1024a_3v1024x8m81_0/bb[0]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[89] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[116]
+ col_1024a_3v1024x8m81_0/WL[21] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[106]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[107] col_1024a_3v1024x8m81_0/saout_R_m2_3v1024x8m81_0/vdd_uq4
+ col_1024a_3v1024x8m81_0/bb[20] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[66]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[125] col_1024a_3v1024x8m81_0/bb[2]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/bb[24] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[84]
+ col_1024a_3v1024x8m81_0/b[9] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[102]
+ col_1024a_3v1024x8m81_0/b[21] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[119]
+ col_1024a_3v1024x8m81_0/bb[4] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[78]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[120] col_1024a_3v1024x8m81_0/WL[8]
+ col_1024a_3v1024x8m81_0/b[5] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[96]
+ WL[27] col_1024a_3v1024x8m81_0/bb[22] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[87]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[114] col_1024a_3v1024x8m81_0/bb[26]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/b[24] WL[44] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[105]
+ col_1024a_3v1024x8m81_0/bb[1] col_1024a_3v1024x8m81_0/bb[6] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[64]
+ col_1024a_3v1024x8m81_0/b[25] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[123]
+ col_1024a_3v1024x8m81_0/b[23] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/bb[8]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[82] col_1024a_3v1024x8m81_0/b[26]
+ col_1024a_3v1024x8m81_0/b[7] col_1024a_3v1024x8m81_0/bb[9] col_1024a_3v1024x8m81_0/WL[58]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[100] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[117]
+ col_1024a_3v1024x8m81_0/b[27] WL[47] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[122]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[76] col_1024a_3v1024x8m81_0/bb[28]
+ col_1024a_3v1024x8m81_0/WL[6] col_1024a_3v1024x8m81_0/b[28] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[67]
+ col_1024a_3v1024x8m81_0/b[13] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[94]
+ col_1024a_3v1024x8m81_0/bb[3] WL[25] col_1024a_3v1024x8m81_0/VDD_uq2 col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[85]
+ col_1024a_3v1024x8m81_0/b[20] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[112]
+ WL[42] col_1024a_3v1024x8m81_0/b[29] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[103]
+ col_1024a_3v1024x8m81_0/WL[62] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[121]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[79] col_1024a_3v1024x8m81_0/bb[17]
+ WL[9] col_1024a_3v1024x8m81_0/bb[21] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[80]
+ col_1024a_3v1024x8m81_0/VDD_uq4 col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[97]
+ col_1024a_3v1024x8m81_0/bb[18] WL[28] WL[54] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[115]
+ col_1024a_3v1024x8m81_0/b[15] col_1024a_3v1024x8m81_0/bb[5] col_1024a_3v1024x8m81_0/saout_m2_3v1024x8m81_4/GWEN
+ col_1024a_3v1024x8m81_0/WL[47] col_1024a_3v1024x8m81_0/bb[19] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[74]
+ col_1024a_3v1024x8m81_0/b[22] WL[4] col_1024a_3v1024x8m81_0/VDD_uq1 col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[65]
+ col_1024a_3v1024x8m81_0/b[31] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[92]
+ col_1024a_3v1024x8m81_0/GWE col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[99]
+ col_1024a_3v1024x8m81_0/VDD_uq0 WL[23] WEN[1] col_1024a_3v1024x8m81_0/b[6] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[110]
+ WL[40] col_1024a_3v1024x8m81_0/bb[23] col_1024a_3v1024x8m81_0/VDD_uq3 col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[101]
+ WL[57] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[83] col_1024a_3v1024x8m81_0/WL[60]
+ WL[15] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[77] col_1024a_3v1024x8m81_0/b[1]
+ col_1024a_3v1024x8m81_0/b[10] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[69]
+ col_1024a_3v1024x8m81_0/bb[7] WL[7] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[95]
+ col_1024a_3v1024x8m81_0/b[2] col_1024a_3v1024x8m81_0/b[11] WL[26] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[113]
+ col_1024a_3v1024x8m81_0/b[3] col_1024a_3v1024x8m81_0/b[12] col_1024a_3v1024x8m81_0/WL[45]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[72] WL[2] VDD col_1024a_3v1024x8m81_0/WL[19]
+ WL[61] VSUBS col_1024a_3v1024x8m81_0/b[4] col_1024a_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[0] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[1] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[2] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[3] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[4] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[5] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[6] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[7] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[8] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[9] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[10] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[11] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[12] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[13] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[14] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[15] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[16] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[17] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[18] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[19] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[20] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[21] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[22] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[23] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[24] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[25] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[26] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[27] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[28] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[29] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[30] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[31] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[32] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[33] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[34] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xdcap_103_novia_3v1024x8m81_0[35] VDD VSUBS VDD dcap_103_novia_3v1024x8m81
Xldummy_3v512x4_3v1024x8m81_0 col_1024a_3v1024x8m81_0/bb[30] VDD col_1024a_3v1024x8m81_0/b[30]
+ WL[4] col_1024a_3v1024x8m81_0/WL[45] VSUBS VSUBS col_1024a_3v1024x8m81_0/b[27] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[117]
+ col_1024a_3v1024x8m81_0/bb[27] VSUBS VDD VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[70]
+ VDD VDD col_1024a_3v1024x8m81_0/WL[62] VDD VSUBS VSUBS col_1024a_3v1024x8m81_0/WL[127]
+ VDD VSUBS col_1024a_3v1024x8m81_0/bb[12] col_1024a_3v1024x8m81_0/bb[0] VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[80]
+ col_1024a_3v1024x8m81_0/b[12] col_1024a_3v1024x8m81_0/b[0] WL[40] VDD VDD VSUBS
+ VSUBS VDD col_1024a_3v1024x8m81_0/b[1] col_1024a_3v1024x8m81_0/bb[1] col_1024a_3v1024x8m81_0/bb[18]
+ col_1024a_3v1024x8m81_0/WL[17] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[90]
+ WL[21] col_1024a_3v1024x8m81_0/b[18] WL[24] VSUBS VSUBS VSUBS VSUBS col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[106]
+ VSUBS col_1024a_3v1024x8m81_0/b[15] WL[0] col_1024a_3v1024x8m81_0/WL[47] col_1024a_3v1024x8m81_0/bb[15]
+ VSUBS VDD VSUBS col_1024a_3v1024x8m81_0/b[29] col_1024a_3v1024x8m81_0/b[11] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[116]
+ VSUBS col_1024a_3v1024x8m81_0/bb[29] col_1024a_3v1024x8m81_0/bb[11] VDD VDD VDD
+ VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[73] VDD col_1024a_3v1024x8m81_0/WL[60]
+ col_1024a_3v1024x8m81_0/bb[22] VSUBS VSUBS col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[126]
+ col_1024a_3v1024x8m81_0/b[22] VDD VSUBS col_1024a_3v1024x8m81_0/bb[14] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/bb[8]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[83] col_1024a_3v1024x8m81_0/b[14]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/b[8] col_1024a_3v1024x8m81_0/WL[40]
+ VDD VDD VSUBS VDD VSUBS col_1024a_3v1024x8m81_0/bb[0] col_1024a_3v1024x8m81_0/b[17]
+ col_1024a_3v1024x8m81_0/b[0] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[93]
+ VDD WL[26] WL[19] col_1024a_3v1024x8m81_0/bb[17] VSUBS VSUBS VSUBS VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[109]
+ VSUBS WL[2] VDD WL[47] VSUBS VSUBS col_1024a_3v1024x8m81_0/bb[28] col_1024a_3v1024x8m81_0/b[13]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[119] VSUBS col_1024a_3v1024x8m81_0/b[28]
+ col_1024a_3v1024x8m81_0/bb[13] VDD VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[72]
+ col_1024a_3v1024x8m81_0/WL[58] col_1024a_3v1024x8m81_0/bb[20] VSUBS VSUBS VDD col_1024a_3v1024x8m81_0/b[20]
+ col_1024a_3v1024x8m81_0/b[9] col_1024a_3v1024x8m81_0/b[7] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[82]
+ col_1024a_3v1024x8m81_0/bb[7] VDD VDD col_1024a_3v1024x8m81_0/WL[38] col_1024a_3v1024x8m81_0/bb[9]
+ VSUBS VSUBS VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/bb[8] VSUBS
+ VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/b[8] col_1024a_3v1024x8m81_0/bb[16]
+ WL[30] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[92] WL[17] col_1024a_3v1024x8m81_0/b[16]
+ VSUBS WL[28] VSUBS VSUBS VDD VSUBS col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[108]
+ VSUBS WL[49] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[65] VSUBS col_1024a_3v1024x8m81_0/bb[30]
+ VSUBS col_1024a_3v1024x8m81_0/bb[12] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[118]
+ VSUBS col_1024a_3v1024x8m81_0/b[30] col_1024a_3v1024x8m81_0/b[12] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[75]
+ WL[54] VDD VSUBS col_1024a_3v1024x8m81_0/b[21] VSUBS col_1024a_3v1024x8m81_0/bb[21]
+ col_1024a_3v1024x8m81_0/bb[6] col_1024a_3v1024x8m81_0/bb[10] col_1024a_3v1024x8m81_0/b[6]
+ VDD col_1024a_3v1024x8m81_0/WL[36] col_1024a_3v1024x8m81_0/b[10] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[85]
+ VDD VSUBS VDD VSUBS VDD col_1024a_3v1024x8m81_0/b[9] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/bb[24]
+ col_1024a_3v1024x8m81_0/bb[9] VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[95]
+ VDD WL[61] WL[34] WL[15] VSUBS col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/b[24]
+ VSUBS VSUBS VSUBS VDD VDD VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[64]
+ VDD WL[51] col_1024a_3v1024x8m81_0/b[31] VDD VSUBS VSUBS col_1024a_3v1024x8m81_0/bb[14]
+ col_1024a_3v1024x8m81_0/bb[31] col_1024a_3v1024x8m81_0/b[14] VDD VDD VDD VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[74]
+ WL[52] VSUBS VDD col_1024a_3v1024x8m81_0/b[19] VSUBS col_1024a_3v1024x8m81_0/bb[19]
+ col_1024a_3v1024x8m81_0/bb[4] col_1024a_3v1024x8m81_0/b[31] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[84]
+ col_1024a_3v1024x8m81_0/b[4] VDD col_1024a_3v1024x8m81_0/bb[31] VDD col_1024a_3v1024x8m81_0/WL[32]
+ VSUBS VDD col_1024a_3v1024x8m81_0/bb[10] col_1024a_3v1024x8m81_0/b[25] col_1024a_3v1024x8m81_0/b[10]
+ WL[1] col_1024a_3v1024x8m81_0/WL[14] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[94]
+ col_1024a_3v1024x8m81_0/bb[25] VSUBS WL[32] VSUBS VSUBS col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[101]
+ VDD VDD VSUBS col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[67] WL[53]
+ VSUBS col_1024a_3v1024x8m81_0/b[23] VSUBS col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[111]
+ col_1024a_3v1024x8m81_0/b[15] VSUBS col_1024a_3v1024x8m81_0/bb[23] col_1024a_3v1024x8m81_0/bb[15]
+ VDD VDD VDD VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[77] VDD WL[50]
+ col_1024a_3v1024x8m81_0/bb[18] VSUBS VSUBS col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[121]
+ VDD col_1024a_3v1024x8m81_0/b[18] VSUBS col_1024a_3v1024x8m81_0/b[5] col_1024a_3v1024x8m81_0/b[23]
+ VDD col_1024a_3v1024x8m81_0/WL[34] VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[87]
+ col_1024a_3v1024x8m81_0/bb[5] col_1024a_3v1024x8m81_0/bb[23] VDD VSUBS VSUBS VDD
+ col_1024a_3v1024x8m81_0/bb[26] WL[5] VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[97]
+ VSUBS col_1024a_3v1024x8m81_0/b[26] col_1024a_3v1024x8m81_0/WL[12] WL[36] VSUBS
+ VSUBS VSUBS VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[100] VDD
+ VSUBS VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[66] VDD WL[55]
+ VSUBS VSUBS col_1024a_3v1024x8m81_0/b[7] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[110]
+ VSUBS col_1024a_3v1024x8m81_0/bb[7] VDD VDD VDD VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[76]
+ WL[48] VDD VSUBS col_1024a_3v1024x8m81_0/b[17] VSUBS col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[120]
+ col_1024a_3v1024x8m81_0/bb[17] VSUBS VDD col_1024a_3v1024x8m81_0/b[3] col_1024a_3v1024x8m81_0/bb[22]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[86] col_1024a_3v1024x8m81_0/bb[3]
+ VDD WL[29] col_1024a_3v1024x8m81_0/b[22] VDD VSUBS VSUBS col_1024a_3v1024x8m81_0/bb[6]
+ col_1024a_3v1024x8m81_0/b[27] col_1024a_3v1024x8m81_0/b[6] VDD WL[7] col_1024a_3v1024x8m81_0/WL[10]
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[96] VSUBS col_1024a_3v1024x8m81_0/bb[27]
+ col_1024a_3v1024x8m81_0/WL[39] VSUBS VSUBS VSUBS VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[103]
+ VDD VSUBS col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[69] VDD WL[57]
+ VSUBS VSUBS col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[113] VSUBS VDD
+ VDD VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[79] VDD WL[46] col_1024a_3v1024x8m81_0/bb[16]
+ VSUBS VSUBS VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[123] VSUBS
+ col_1024a_3v1024x8m81_0/b[16] col_1024a_3v1024x8m81_0/bb[20] col_1024a_3v1024x8m81_0/bb[2]
+ col_1024a_3v1024x8m81_0/b[2] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[89]
+ VDD VDD WL[27] col_1024a_3v1024x8m81_0/b[20] VSUBS VSUBS VDD col_1024a_3v1024x8m81_0/bb[4]
+ col_1024a_3v1024x8m81_0/b[4] col_1024a_3v1024x8m81_0/b[29] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[99]
+ WL[9] col_1024a_3v1024x8m81_0/WL[8] col_1024a_3v1024x8m81_0/bb[29] VDD VSUBS VSUBS
+ VSUBS VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[102] VSUBS VDD
+ col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[68] VDD VSUBS col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[112]
+ VSUBS VDD VDD VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[78] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/bb[24]
+ VSUBS col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[122] VSUBS col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/b[24]
+ col_1024a_3v1024x8m81_0/b[21] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[88]
+ col_1024a_3v1024x8m81_0/bb[21] VSUBS col_1024a_3v1024x8m81_0/b[5] col_1024a_3v1024x8m81_0/bb[5]
+ col_1024a_3v1024x8m81_0/bb[28] WL[11] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[98]
+ VSUBS col_1024a_3v1024x8m81_0/WL[19] col_1024a_3v1024x8m81_0/b[28] VSUBS VSUBS col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[105]
+ VDD VSUBS col_1024a_3v1024x8m81_0/WL[41] VSUBS VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[115]
+ VSUBS VDD VDD VDD VDD WL[59] VDD col_1024a_3v1024x8m81_0/b[25] VSUBS VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[125]
+ VSUBS col_1024a_3v1024x8m81_0/bb[25] VDD col_1024a_3v1024x8m81_0/b[11] col_1024a_3v1024x8m81_0/bb[11]
+ WL[44] VDD VDD VDD VDD VSUBS VDD col_1024a_3v1024x8m81_0/b[3] col_1024a_3v1024x8m81_0/bb[3]
+ VSUBS VDD col_1024a_3v1024x8m81_0/WL[13] VDD WL[25] col_1024a_3v1024x8m81_0/WL[21]
+ VSUBS VSUBS VSUBS VDD VDD VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[104]
+ VSUBS col_1024a_3v1024x8m81_0/WL[6] col_1024a_3v1024x8m81_0/WL[43] VSUBS VSUBS col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[114]
+ VSUBS VDD VDD VDD VDD WL[3] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[71]
+ VDD VSUBS VSUBS col_1024a_3v1024x8m81_0/bb[26] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[124]
+ col_1024a_3v1024x8m81_0/b[26] VSUBS col_1024a_3v1024x8m81_0/b[13] VDD col_1024a_3v1024x8m81_0/b[1]
+ VSUBS col_1024a_3v1024x8m81_0/bb[13] col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[81]
+ VDD col_1024a_3v1024x8m81_0/bb[1] VDD WL[42] VDD VSUBS VDD VSUBS col_1024a_3v1024x8m81_0/bb[2]
+ col_1024a_3v1024x8m81_0/b[19] col_1024a_3v1024x8m81_0/b[2] col_1024a_3v1024x8m81_0/WL[15]
+ WL[23] VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[91] VSUBS VSUBS
+ col_1024a_3v1024x8m81_0/bb[19] VDD WL[22] VSUBS VSUBS VDD col_1024a_3v1024x8m81_0/Cell_array8x8_3v1024x8m81_0/wl[107]
+ VSUBS VSUBS ldummy_3v512x4_3v1024x8m81
.ends

.subckt pmos_5p04310591302072_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.1406p pd=10.61u as=2.1406p ps=10.61u w=4.865u l=0.28u
.ends

.subckt pmos_1p2$$47512620_3v1024x8m81 w_n133_n66# a_n14_n34# pmos_5p04310591302072_3v1024x8m81_0/S
+ pmos_5p04310591302072_3v1024x8m81_0/D
Xpmos_5p04310591302072_3v1024x8m81_0 pmos_5p04310591302072_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302072_3v1024x8m81_0/S pmos_5p04310591302072_3v1024x8m81
.ends

.subckt pmos_5p04310591302068_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.3276p pd=11.46u as=2.3276p ps=11.46u w=5.29u l=0.28u
.ends

.subckt pmos_1p2$$47513644_3v1024x8m81 pmos_5p04310591302068_3v1024x8m81_0/D a_n14_n34#
+ pmos_5p04310591302068_3v1024x8m81_0/S w_n133_n65#
Xpmos_5p04310591302068_3v1024x8m81_0 pmos_5p04310591302068_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302068_3v1024x8m81_0/S pmos_5p04310591302068_3v1024x8m81
.ends

.subckt nmos_5p04310591302057_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.9306p pd=5.11u as=0.9306p ps=5.11u w=2.115u l=0.28u
.ends

.subckt nmos_1p2$$47514668_3v1024x8m81 nmos_5p04310591302057_3v1024x8m81_0/S nmos_5p04310591302057_3v1024x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p04310591302057_3v1024x8m81_0 nmos_5p04310591302057_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p04310591302057_3v1024x8m81_0/S VSUBS nmos_5p04310591302057_3v1024x8m81
.ends

.subckt xpredec1_xa_3v1024x8m81 m1_n40_n4147# m1_n40_n4005# m3_n46_n5510# a_145_n5643#
+ m1_n40_n3864# m1_n40_n3582# m1_n40_n3723# a_0_56# m1_n40_n3441# M3_M2$$47333420_3v1024x8m81_1/VSUBS
+ a_465_n5643# pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/D
+ pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/S a_305_n5643#
Xpmos_1p2$$47512620_3v1024x8m81_0 pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/S
+ a_145_n5643# pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/S
+ pmos_1p2$$47512620_3v1024x8m81_3/pmos_5p04310591302072_3v1024x8m81_0/S pmos_1p2$$47512620_3v1024x8m81
Xpmos_1p2$$47512620_3v1024x8m81_1 pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/S
+ a_465_n5643# pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/S
+ pmos_1p2$$47512620_3v1024x8m81_3/pmos_5p04310591302072_3v1024x8m81_0/S pmos_1p2$$47512620_3v1024x8m81
Xpmos_1p2$$47512620_3v1024x8m81_3 pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/S
+ a_305_n5643# pmos_1p2$$47512620_3v1024x8m81_3/pmos_5p04310591302072_3v1024x8m81_0/S
+ pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/S pmos_1p2$$47512620_3v1024x8m81
Xpmos_1p2$$47513644_3v1024x8m81_1 pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/D
+ pmos_1p2$$47512620_3v1024x8m81_3/pmos_5p04310591302072_3v1024x8m81_0/S pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/S
+ pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/S pmos_1p2$$47513644_3v1024x8m81
Xpmos_1p2$$47513644_3v1024x8m81_0 pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/S
+ pmos_1p2$$47512620_3v1024x8m81_3/pmos_5p04310591302072_3v1024x8m81_0/S pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/D
+ pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/S pmos_1p2$$47513644_3v1024x8m81
Xpmos_1p2$$47513644_3v1024x8m81_2 pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/D
+ pmos_1p2$$47512620_3v1024x8m81_3/pmos_5p04310591302072_3v1024x8m81_0/S pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/S
+ pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/S pmos_1p2$$47513644_3v1024x8m81
Xnmos_1p2$$47514668_3v1024x8m81_0 M3_M2$$47333420_3v1024x8m81_1/VSUBS pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/D
+ pmos_1p2$$47512620_3v1024x8m81_3/pmos_5p04310591302072_3v1024x8m81_0/S M3_M2$$47333420_3v1024x8m81_1/VSUBS
+ nmos_1p2$$47514668_3v1024x8m81
Xnmos_1p2$$47514668_3v1024x8m81_1 pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/D
+ M3_M2$$47333420_3v1024x8m81_1/VSUBS pmos_1p2$$47512620_3v1024x8m81_3/pmos_5p04310591302072_3v1024x8m81_0/S
+ M3_M2$$47333420_3v1024x8m81_1/VSUBS nmos_1p2$$47514668_3v1024x8m81
Xnmos_1p2$$47514668_3v1024x8m81_2 M3_M2$$47333420_3v1024x8m81_1/VSUBS pmos_1p2$$47513644_3v1024x8m81_2/pmos_5p04310591302068_3v1024x8m81_0/D
+ pmos_1p2$$47512620_3v1024x8m81_3/pmos_5p04310591302072_3v1024x8m81_0/S M3_M2$$47333420_3v1024x8m81_1/VSUBS
+ nmos_1p2$$47514668_3v1024x8m81
X0 a_361_n5592# a_305_n5643# a_201_n5592# M3_M2$$47333420_3v1024x8m81_1/VSUBS nfet_03v3 ad=1.5145p pd=6.345u as=1.5145p ps=6.345u w=5.825u l=0.28u
X1 a_201_n5592# a_145_n5643# M3_M2$$47333420_3v1024x8m81_1/VSUBS M3_M2$$47333420_3v1024x8m81_1/VSUBS nfet_03v3 ad=1.5145p pd=6.345u as=2.65037p ps=12.56u w=5.825u l=0.28u
X2 pmos_1p2$$47512620_3v1024x8m81_3/pmos_5p04310591302072_3v1024x8m81_0/S a_465_n5643# a_361_n5592# M3_M2$$47333420_3v1024x8m81_1/VSUBS nfet_03v3 ad=2.82512p pd=12.62u as=1.5145p ps=6.345u w=5.825u l=0.28u
.ends

.subckt nmos_5p04310591302053_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.2772p pd=2.14u as=0.2772p ps=2.14u w=0.63u l=0.28u
.ends

.subckt nmos_1p2$$47342636_3v1024x8m81 nmos_5p04310591302053_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p04310591302053_3v1024x8m81_0/S VSUBS
Xnmos_5p04310591302053_3v1024x8m81_0 nmos_5p04310591302053_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p04310591302053_3v1024x8m81_0/S VSUBS nmos_5p04310591302053_3v1024x8m81
.ends

.subckt pmos_5p04310591302070_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=3.3528p pd=16.12u as=3.3528p ps=16.12u w=7.62u l=0.28u
.ends

.subckt pmos_1p2$$47337516_3v1024x8m81 pmos_5p04310591302070_3v1024x8m81_0/D a_n14_n34#
+ pmos_5p04310591302070_3v1024x8m81_0/S w_n133_n65#
Xpmos_5p04310591302070_3v1024x8m81_0 pmos_5p04310591302070_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302070_3v1024x8m81_0/S pmos_5p04310591302070_3v1024x8m81
.ends

.subckt nmos_1p2_157_3v1024x8m81 nmos_5p04310591302010_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v1024x8m81_0/S VSUBS
Xnmos_5p04310591302010_3v1024x8m81_0 nmos_5p04310591302010_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v1024x8m81_0/S VSUBS nmos_5p04310591302010_3v1024x8m81
.ends

.subckt pmos_5p04310591302058_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.5499p pd=2.635u as=0.9306p ps=5.11u w=2.115u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.9306p pd=5.11u as=0.5499p ps=2.635u w=2.115u l=0.28u
.ends

.subckt pmos_1p2$$47331372_3v1024x8m81 a_n42_n34# w_n133_n66# pmos_5p04310591302058_3v1024x8m81_0/S
+ pmos_5p04310591302058_3v1024x8m81_0/D a_118_n34# pmos_5p04310591302058_3v1024x8m81_0/S_uq0
Xpmos_5p04310591302058_3v1024x8m81_0 pmos_5p04310591302058_3v1024x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302058_3v1024x8m81_0/S_uq0 pmos_5p04310591302058_3v1024x8m81_0/S
+ pmos_5p04310591302058_3v1024x8m81
.ends

.subckt pmos_1p2_161_3v1024x8m81 pmos_5p04310591302041_3v1024x8m81_0/D a_n14_89# pmos_5p04310591302041_3v1024x8m81_0/S
+ w_n133_n65#
Xpmos_5p04310591302041_3v1024x8m81_0 pmos_5p04310591302041_3v1024x8m81_0/D a_n14_89#
+ w_n133_n65# pmos_5p04310591302041_3v1024x8m81_0/S pmos_5p04310591302041_3v1024x8m81
.ends

.subckt nmos_5p04310591302059_3v1024x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.28u
.ends

.subckt nmos_1p2$$47329324_3v1024x8m81 nmos_5p04310591302059_3v1024x8m81_0/S_uq0 nmos_5p04310591302059_3v1024x8m81_0/D
+ a_118_n34# a_n41_n34# nmos_5p04310591302059_3v1024x8m81_0/S VSUBS
Xnmos_5p04310591302059_3v1024x8m81_0 nmos_5p04310591302059_3v1024x8m81_0/D a_n41_n34#
+ a_118_n34# nmos_5p04310591302059_3v1024x8m81_0/S_uq0 nmos_5p04310591302059_3v1024x8m81_0/S
+ VSUBS nmos_5p04310591302059_3v1024x8m81
.ends

.subckt pmos_1p2_160_3v1024x8m81 w_n133_n66# pmos_5p04310591302014_3v1024x8m81_0/S
+ a_n14_n34# pmos_5p04310591302014_3v1024x8m81_0/D
Xpmos_5p04310591302014_3v1024x8m81_0 pmos_5p04310591302014_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302014_3v1024x8m81_0/S pmos_5p04310591302014_3v1024x8m81
.ends

.subckt alatch_3v1024x8m81 en ab a vdd enb a_886_665# vss
Xnmos_1p2_157_3v1024x8m81_0 a a_886_665# nmos_5p0431059130208_3v1024x8m81_1/S vss
+ nmos_1p2_157_3v1024x8m81
Xnmos_5p0431059130208_3v1024x8m81_0 vss ab nmos_5p0431059130208_3v1024x8m81_1/D vss
+ nmos_5p0431059130208_3v1024x8m81
Xnmos_5p0431059130208_3v1024x8m81_1 nmos_5p0431059130208_3v1024x8m81_1/D enb nmos_5p0431059130208_3v1024x8m81_1/S
+ vss nmos_5p0431059130208_3v1024x8m81
Xpmos_1p2$$47331372_3v1024x8m81_0 nmos_5p0431059130208_3v1024x8m81_1/S vdd vdd ab
+ nmos_5p0431059130208_3v1024x8m81_1/S vdd pmos_1p2$$47331372_3v1024x8m81
Xpmos_1p2_161_3v1024x8m81_0 nmos_5p0431059130208_3v1024x8m81_1/D a_886_665# nmos_5p0431059130208_3v1024x8m81_1/S
+ vdd pmos_1p2_161_3v1024x8m81
Xpmos_1p2_161_3v1024x8m81_1 vdd ab nmos_5p0431059130208_3v1024x8m81_1/D vdd pmos_1p2_161_3v1024x8m81
Xnmos_1p2$$47329324_3v1024x8m81_0 vss ab nmos_5p0431059130208_3v1024x8m81_1/S nmos_5p0431059130208_3v1024x8m81_1/S
+ vss vss nmos_1p2$$47329324_3v1024x8m81
Xpmos_1p2_160_3v1024x8m81_0 vdd nmos_5p0431059130208_3v1024x8m81_1/S enb a pmos_1p2_160_3v1024x8m81
.ends

.subckt nmos_5p04310591302071_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.3508p pd=7.02u as=1.3508p ps=7.02u w=3.07u l=0.28u
.ends

.subckt nmos_1p2$$47336492_3v1024x8m81 nmos_5p04310591302071_3v1024x8m81_0/S a_n14_n34#
+ nmos_5p04310591302071_3v1024x8m81_0/D VSUBS
Xnmos_5p04310591302071_3v1024x8m81_0 nmos_5p04310591302071_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p04310591302071_3v1024x8m81_0/S VSUBS nmos_5p04310591302071_3v1024x8m81
.ends

.subckt xpredec1_bot_3v1024x8m81 m1_n74_2740# alatch_3v1024x8m81_0/a pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/S
+ m1_n74_3446# alatch_3v1024x8m81_0/enb m1_n74_3164# alatch_3v1024x8m81_0/vdd m1_n74_3305#
+ pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D m1_n74_3023#
+ VSUBS m3_9_2964# m1_n74_2881# pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
Xpmos_1p2$$47337516_3v1024x8m81_0 pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/S
+ pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/S pmos_1p2$$47337516_3v1024x8m81
Xpmos_1p2$$47337516_3v1024x8m81_1 pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ alatch_3v1024x8m81_0/ab pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/S
+ pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/S pmos_1p2$$47337516_3v1024x8m81
Xalatch_3v1024x8m81_0 alatch_3v1024x8m81_0/en alatch_3v1024x8m81_0/ab alatch_3v1024x8m81_0/a
+ alatch_3v1024x8m81_0/vdd alatch_3v1024x8m81_0/enb m3_9_2964# VSUBS alatch_3v1024x8m81
Xnmos_1p2$$47336492_3v1024x8m81_0 VSUBS pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D VSUBS nmos_1p2$$47336492_3v1024x8m81
Xnmos_1p2$$47336492_3v1024x8m81_1 VSUBS alatch_3v1024x8m81_0/ab pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ VSUBS nmos_1p2$$47336492_3v1024x8m81
.ends

.subckt nmos_5p04310591302056_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.3916p pd=2.66u as=0.3916p ps=2.66u w=0.89u l=0.28u
.ends

.subckt pmos_5p04310591302062_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.2067p pd=1.315u as=0.3498p ps=2.47u w=0.795u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.3498p pd=2.47u as=0.2067p ps=1.315u w=0.795u l=0.28u
.ends

.subckt pmos_1p2$$47109164_3v1024x8m81 pmos_5p04310591302062_3v1024x8m81_0/w_n202_n86#
+ pmos_5p04310591302062_3v1024x8m81_0/D pmos_5p04310591302062_3v1024x8m81_0/S_uq0
+ a_118_159# pmos_5p04310591302062_3v1024x8m81_0/S a_n42_159#
Xpmos_5p04310591302062_3v1024x8m81_0 pmos_5p04310591302062_3v1024x8m81_0/D a_n42_159#
+ a_118_159# pmos_5p04310591302062_3v1024x8m81_0/w_n202_n86# pmos_5p04310591302062_3v1024x8m81_0/S_uq0
+ pmos_5p04310591302062_3v1024x8m81_0/S pmos_5p04310591302062_3v1024x8m81
.ends

.subckt xpredec1_3v1024x8m81 men x[7] x[6] x[5] x[4] x[3] x[2] x[1] x[0] clk vdd_uq0
+ w_5024_6624# A[0] A[1] vdd xpredec1_xa_3v1024x8m81_7/m3_n46_n5510# A[2] vss xpredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/vdd
+ pmos_1p2$$47109164_3v1024x8m81_0/pmos_5p04310591302062_3v1024x8m81_0/w_n202_n86#
Xxpredec1_xa_3v1024x8m81_2 xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81_7/m3_n46_n5510# xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ vss xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ vss xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ x[5] vdd_uq0 xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81
Xxpredec1_xa_3v1024x8m81_3 xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81_7/m3_n46_n5510# xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81_3/a_0_56# xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ vss xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ x[7] vdd_uq0 xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81
Xnmos_1p2$$47342636_3v1024x8m81_0 vss nmos_5p04310591302056_3v1024x8m81_1/D xpredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/enb
+ vss nmos_1p2$$47342636_3v1024x8m81
Xxpredec1_xa_3v1024x8m81_4 xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81_7/m3_n46_n5510# xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81_4/a_0_56# xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ vss xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ x[2] vdd_uq0 xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81
Xxpredec1_xa_3v1024x8m81_5 xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81_7/m3_n46_n5510# xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81_5/a_0_56# xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ vss xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ x[0] vdd_uq0 xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81
Xxpredec1_xa_3v1024x8m81_6 xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81_7/m3_n46_n5510# xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81_6/a_0_56# xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ vss xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ x[4] vdd_uq0 xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81
Xxpredec1_xa_3v1024x8m81_7 xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81_7/m3_n46_n5510# xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81_7/a_0_56# xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ vss xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ x[6] vdd_uq0 xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81
Xxpredec1_bot_3v1024x8m81_0 xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ A[0] vdd_uq0 xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/enb xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/vdd xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ vss nmos_5p04310591302056_3v1024x8m81_1/D xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81
Xxpredec1_bot_3v1024x8m81_1 xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ A[2] vdd_uq0 xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/enb xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/vdd xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ vss nmos_5p04310591302056_3v1024x8m81_1/D xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81
Xxpredec1_bot_3v1024x8m81_2 xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ A[1] vdd_uq0 xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/enb xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/vdd xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ vss nmos_5p04310591302056_3v1024x8m81_1/D xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81
Xnmos_5p04310591302056_3v1024x8m81_0 vss clk nmos_5p04310591302056_3v1024x8m81_1/D
+ vss nmos_5p04310591302056_3v1024x8m81
Xnmos_5p04310591302056_3v1024x8m81_1 nmos_5p04310591302056_3v1024x8m81_1/D men vss
+ vss nmos_5p04310591302056_3v1024x8m81
Xpmos_1p2$$47109164_3v1024x8m81_0 pmos_1p2$$47109164_3v1024x8m81_0/pmos_5p04310591302062_3v1024x8m81_0/w_n202_n86#
+ xpredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/enb vdd nmos_5p04310591302056_3v1024x8m81_1/D
+ vdd nmos_5p04310591302056_3v1024x8m81_1/D pmos_1p2$$47109164_3v1024x8m81
Xxpredec1_xa_3v1024x8m81_0 xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81_7/m3_n46_n5510# xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81_0/a_0_56# xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ vss xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ x[3] vdd_uq0 xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81
Xxpredec1_xa_3v1024x8m81_1 xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81_7/m3_n46_n5510# xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_bot_3v1024x8m81_0/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ vss xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_1/pmos_5p04310591302070_3v1024x8m81_0/D
+ vss xpredec1_bot_3v1024x8m81_1/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ x[1] vdd_uq0 xpredec1_bot_3v1024x8m81_2/pmos_1p2$$47337516_3v1024x8m81_0/pmos_5p04310591302070_3v1024x8m81_0/D
+ xpredec1_xa_3v1024x8m81
X0 a_5287_6723# men vdd w_5024_6624# pfet_03v3 ad=0.212p pd=1.46u as=0.5936p ps=3.24u w=1.06u l=0.28u
X1 a_5600_6723# clk nmos_5p04310591302056_3v1024x8m81_1/D w_5024_6624# pfet_03v3 ad=0.19345p pd=1.425u as=0.32065p ps=1.665u w=1.06u l=0.28u
X2 nmos_5p04310591302056_3v1024x8m81_1/D clk a_5287_6723# w_5024_6624# pfet_03v3 ad=0.32065p pd=1.665u as=0.212p ps=1.46u w=1.06u l=0.28u
X3 vdd men a_5600_6723# w_5024_6624# pfet_03v3 ad=0.5883p pd=3.23u as=0.19345p ps=1.425u w=1.06u l=0.28u
.ends

.subckt pmos_5p04310591302069_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.1378p pd=1.05u as=0.2332p ps=1.94u w=0.53u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.2332p pd=1.94u as=0.1378p ps=1.05u w=0.53u l=0.28u
.ends

.subckt pmos_5p04310591302067_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=3.1196p pd=15.06u as=3.1196p ps=15.06u w=7.09u l=0.28u
.ends

.subckt pmos_1p2$$47643692_3v1024x8m81 w_n133_n66# pmos_5p04310591302067_3v1024x8m81_0/D
+ a_n14_n34# pmos_5p04310591302067_3v1024x8m81_0/S
Xpmos_5p04310591302067_3v1024x8m81_0 pmos_5p04310591302067_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302067_3v1024x8m81_0/S pmos_5p04310591302067_3v1024x8m81
.ends

.subckt pmos_1p2$$47642668_3v1024x8m81 pmos_5p04310591302067_3v1024x8m81_0/D a_n14_n34#
+ w_n194_n66# pmos_5p04310591302067_3v1024x8m81_0/S
Xpmos_5p04310591302067_3v1024x8m81_0 pmos_5p04310591302067_3v1024x8m81_0/D a_n14_n34#
+ w_n194_n66# pmos_5p04310591302067_3v1024x8m81_0/S pmos_5p04310591302067_3v1024x8m81
.ends

.subckt nmos_1p2$$47641644_3v1024x8m81 nmos_5p04310591302057_3v1024x8m81_0/S nmos_5p04310591302057_3v1024x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p04310591302057_3v1024x8m81_0 nmos_5p04310591302057_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p04310591302057_3v1024x8m81_0/S VSUBS nmos_5p04310591302057_3v1024x8m81
.ends

.subckt xpredec0_xa_3v1024x8m81 m3_107_5938# m1_255_3759# a_612_1974# m1_255_3263#
+ m1_255_3619# m1_255_3901# m3_598_2319# a_472_3898# M3_M2$$47644716_3v1024x8m81_2/VSUBS
+ pmos_1p2$$47513644_3v1024x8m81_3/pmos_5p04310591302068_3v1024x8m81_0/D pmos_1p2$$47513644_3v1024x8m81_3/pmos_5p04310591302068_3v1024x8m81_0/S
+ pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/D nmos_1p2$$47641644_3v1024x8m81_3/nmos_5p04310591302057_3v1024x8m81_0/D
Xpmos_1p2$$47643692_3v1024x8m81_0 pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/D
+ pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/D a_472_3898#
+ pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/S pmos_1p2$$47643692_3v1024x8m81
Xpmos_1p2$$47642668_3v1024x8m81_0 pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/S
+ a_612_1974# pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/D
+ pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/D pmos_1p2$$47642668_3v1024x8m81
Xpmos_1p2$$47513644_3v1024x8m81_0 pmos_1p2$$47513644_3v1024x8m81_3/pmos_5p04310591302068_3v1024x8m81_0/S
+ pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/S pmos_1p2$$47513644_3v1024x8m81_3/pmos_5p04310591302068_3v1024x8m81_0/D
+ pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/D pmos_1p2$$47513644_3v1024x8m81
Xpmos_1p2$$47513644_3v1024x8m81_1 pmos_1p2$$47513644_3v1024x8m81_3/pmos_5p04310591302068_3v1024x8m81_0/D
+ pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/S pmos_1p2$$47513644_3v1024x8m81_3/pmos_5p04310591302068_3v1024x8m81_0/S
+ pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/D pmos_1p2$$47513644_3v1024x8m81
Xpmos_1p2$$47513644_3v1024x8m81_2 pmos_1p2$$47513644_3v1024x8m81_3/pmos_5p04310591302068_3v1024x8m81_0/S
+ pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/S pmos_1p2$$47513644_3v1024x8m81_3/pmos_5p04310591302068_3v1024x8m81_0/D
+ pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/D pmos_1p2$$47513644_3v1024x8m81
Xpmos_1p2$$47513644_3v1024x8m81_3 pmos_1p2$$47513644_3v1024x8m81_3/pmos_5p04310591302068_3v1024x8m81_0/D
+ pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/S pmos_1p2$$47513644_3v1024x8m81_3/pmos_5p04310591302068_3v1024x8m81_0/S
+ pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/D pmos_1p2$$47513644_3v1024x8m81
Xnmos_1p2$$47641644_3v1024x8m81_0 nmos_1p2$$47641644_3v1024x8m81_3/nmos_5p04310591302057_3v1024x8m81_0/D
+ pmos_1p2$$47513644_3v1024x8m81_3/pmos_5p04310591302068_3v1024x8m81_0/D pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/S
+ M3_M2$$47644716_3v1024x8m81_2/VSUBS nmos_1p2$$47641644_3v1024x8m81
Xnmos_1p2$$47641644_3v1024x8m81_1 nmos_1p2$$47641644_3v1024x8m81_3/nmos_5p04310591302057_3v1024x8m81_0/D
+ pmos_1p2$$47513644_3v1024x8m81_3/pmos_5p04310591302068_3v1024x8m81_0/D pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/S
+ M3_M2$$47644716_3v1024x8m81_2/VSUBS nmos_1p2$$47641644_3v1024x8m81
Xnmos_1p2$$47641644_3v1024x8m81_2 pmos_1p2$$47513644_3v1024x8m81_3/pmos_5p04310591302068_3v1024x8m81_0/D
+ nmos_1p2$$47641644_3v1024x8m81_3/nmos_5p04310591302057_3v1024x8m81_0/D pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/S
+ M3_M2$$47644716_3v1024x8m81_2/VSUBS nmos_1p2$$47641644_3v1024x8m81
Xnmos_1p2$$47641644_3v1024x8m81_3 pmos_1p2$$47513644_3v1024x8m81_3/pmos_5p04310591302068_3v1024x8m81_0/D
+ nmos_1p2$$47641644_3v1024x8m81_3/nmos_5p04310591302057_3v1024x8m81_0/D pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/S
+ M3_M2$$47644716_3v1024x8m81_2/VSUBS nmos_1p2$$47641644_3v1024x8m81
X0 M3_M2$$47644716_3v1024x8m81_2/VSUBS a_612_1974# a_539_2025# M3_M2$$47644716_3v1024x8m81_2/VSUBS nfet_03v3 ad=3.1746p pd=12.55u as=1.0439p ps=6.085u w=5.72u l=0.28u
X1 a_539_2025# a_472_3898# pmos_1p2$$47643692_3v1024x8m81_0/pmos_5p04310591302067_3v1024x8m81_0/S M3_M2$$47644716_3v1024x8m81_2/VSUBS nfet_03v3 ad=1.0439p pd=6.085u as=3.146p ps=12.54u w=5.72u l=0.28u
.ends

.subckt nmos_5p04310591302066_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.4454p pd=7.45u as=1.4454p ps=7.45u w=3.285u l=0.28u
.ends

.subckt pmos_5p04310591302063_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.7016p pd=13.16u as=2.7016p ps=13.16u w=6.14u l=0.28u
.ends

.subckt pmos_1p2$$47504428_3v1024x8m81 pmos_5p04310591302063_3v1024x8m81_0/D w_n133_n66#
+ a_n14_n34# pmos_5p04310591302063_3v1024x8m81_0/S
Xpmos_5p04310591302063_3v1024x8m81_0 pmos_5p04310591302063_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302063_3v1024x8m81_0/S pmos_5p04310591302063_3v1024x8m81
.ends

.subckt nmos_5p04310591302065_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.0714p pd=5.75u as=1.0714p ps=5.75u w=2.435u l=0.28u
.ends

.subckt nmos_1p2$$47502380_3v1024x8m81 nmos_5p04310591302065_3v1024x8m81_0/S nmos_5p04310591302065_3v1024x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p04310591302065_3v1024x8m81_0 nmos_5p04310591302065_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p04310591302065_3v1024x8m81_0/S VSUBS nmos_5p04310591302065_3v1024x8m81
.ends

.subckt pmos_5p04310591302064_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=3.6322p pd=17.39u as=3.6322p ps=17.39u w=8.255u l=0.28u
.ends

.subckt pmos_1p2$$47503404_3v1024x8m81 a_n14_n34# pmos_5p04310591302064_3v1024x8m81_0/S
+ pmos_5p04310591302064_3v1024x8m81_0/D w_n133_n65#
Xpmos_5p04310591302064_3v1024x8m81_0 pmos_5p04310591302064_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302064_3v1024x8m81_0/S pmos_5p04310591302064_3v1024x8m81
.ends

.subckt xpredec0_bot_3v1024x8m81 nmos_1p2$$47502380_3v1024x8m81_0/nmos_5p04310591302065_3v1024x8m81_0/S
+ nmos_5p04310591302066_3v1024x8m81_0/D m1_n74_3354# m1_n74_3071# alatch_3v1024x8m81_0/a
+ pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/S m1_n74_3213#
+ m1_n74_2930# pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ m3_10_3351# alatch_3v1024x8m81_0/enb alatch_3v1024x8m81_0/vdd pmos_1p2$$47503404_3v1024x8m81_0/pmos_5p04310591302064_3v1024x8m81_0/S
+ VSUBS
Xnmos_5p04310591302066_3v1024x8m81_0 nmos_5p04310591302066_3v1024x8m81_0/D alatch_3v1024x8m81_0/ab
+ VSUBS VSUBS nmos_5p04310591302066_3v1024x8m81
Xpmos_1p2$$47504428_3v1024x8m81_0 pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ pmos_1p2$$47503404_3v1024x8m81_0/pmos_5p04310591302064_3v1024x8m81_0/S nmos_5p04310591302066_3v1024x8m81_0/D
+ pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/S pmos_1p2$$47504428_3v1024x8m81
Xnmos_1p2$$47502380_3v1024x8m81_0 nmos_1p2$$47502380_3v1024x8m81_0/nmos_5p04310591302065_3v1024x8m81_0/S
+ pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D nmos_5p04310591302066_3v1024x8m81_0/D
+ VSUBS nmos_1p2$$47502380_3v1024x8m81
Xalatch_3v1024x8m81_0 alatch_3v1024x8m81_0/en alatch_3v1024x8m81_0/ab alatch_3v1024x8m81_0/a
+ alatch_3v1024x8m81_0/vdd alatch_3v1024x8m81_0/enb m3_10_3351# VSUBS alatch_3v1024x8m81
Xpmos_1p2$$47503404_3v1024x8m81_0 alatch_3v1024x8m81_0/ab pmos_1p2$$47503404_3v1024x8m81_0/pmos_5p04310591302064_3v1024x8m81_0/S
+ nmos_5p04310591302066_3v1024x8m81_0/D pmos_1p2$$47503404_3v1024x8m81_0/pmos_5p04310591302064_3v1024x8m81_0/S
+ pmos_1p2$$47503404_3v1024x8m81
.ends

.subckt xpredec0_3v1024x8m81 vss A[0] x[1] x[2] x[3] A[1] clk vss_uq0 vdd_uq0 vdd_uq2
+ x[0] men vdd VSUBS
Xnmos_5p04310591302040_3v1024x8m81_1 VSUBS clk nmos_5p04310591302040_3v1024x8m81_1/S
+ VSUBS nmos_5p04310591302040_3v1024x8m81
Xnmos_5p04310591302040_3v1024x8m81_0 nmos_5p04310591302040_3v1024x8m81_1/S men VSUBS
+ VSUBS nmos_5p04310591302040_3v1024x8m81
Xpmos_5p04310591302069_3v1024x8m81_0 pmos_5p04310591302069_3v1024x8m81_0/D nmos_5p04310591302040_3v1024x8m81_1/S
+ nmos_5p04310591302040_3v1024x8m81_1/S vdd_uq2 vdd_uq2 vdd_uq2 pmos_5p04310591302069_3v1024x8m81
Xxpredec0_xa_3v1024x8m81_0 VSUBS xpredec0_bot_3v1024x8m81_1/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ xpredec0_bot_3v1024x8m81_0/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ xpredec0_bot_3v1024x8m81_0/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ xpredec0_bot_3v1024x8m81_0/nmos_5p04310591302066_3v1024x8m81_0/D xpredec0_bot_3v1024x8m81_1/nmos_5p04310591302066_3v1024x8m81_0/D
+ vdd xpredec0_bot_3v1024x8m81_1/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ VSUBS x[0] vdd_uq2 vdd_uq2 VSUBS xpredec0_xa_3v1024x8m81
Xxpredec0_xa_3v1024x8m81_1 VSUBS xpredec0_bot_3v1024x8m81_1/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ xpredec0_bot_3v1024x8m81_0/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ xpredec0_bot_3v1024x8m81_0/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ xpredec0_bot_3v1024x8m81_0/nmos_5p04310591302066_3v1024x8m81_0/D xpredec0_bot_3v1024x8m81_1/nmos_5p04310591302066_3v1024x8m81_0/D
+ vdd xpredec0_bot_3v1024x8m81_1/nmos_5p04310591302066_3v1024x8m81_0/D VSUBS x[2]
+ vdd_uq2 vdd_uq2 VSUBS xpredec0_xa_3v1024x8m81
Xxpredec0_xa_3v1024x8m81_2 VSUBS xpredec0_bot_3v1024x8m81_1/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ xpredec0_bot_3v1024x8m81_0/nmos_5p04310591302066_3v1024x8m81_0/D xpredec0_bot_3v1024x8m81_0/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ xpredec0_bot_3v1024x8m81_0/nmos_5p04310591302066_3v1024x8m81_0/D xpredec0_bot_3v1024x8m81_1/nmos_5p04310591302066_3v1024x8m81_0/D
+ vdd xpredec0_bot_3v1024x8m81_1/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ VSUBS x[1] vdd_uq2 vdd_uq2 VSUBS xpredec0_xa_3v1024x8m81
Xnmos_1p2$$46563372_3v1024x8m81_0 pmos_5p04310591302069_3v1024x8m81_0/D VSUBS nmos_5p04310591302040_3v1024x8m81_1/S
+ VSUBS nmos_1p2$$46563372_3v1024x8m81
Xxpredec0_xa_3v1024x8m81_3 VSUBS xpredec0_bot_3v1024x8m81_1/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ xpredec0_bot_3v1024x8m81_0/nmos_5p04310591302066_3v1024x8m81_0/D xpredec0_bot_3v1024x8m81_0/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ xpredec0_bot_3v1024x8m81_0/nmos_5p04310591302066_3v1024x8m81_0/D xpredec0_bot_3v1024x8m81_1/nmos_5p04310591302066_3v1024x8m81_0/D
+ vdd xpredec0_bot_3v1024x8m81_1/nmos_5p04310591302066_3v1024x8m81_0/D VSUBS x[3]
+ vdd_uq2 vdd_uq2 VSUBS xpredec0_xa_3v1024x8m81
Xxpredec0_bot_3v1024x8m81_0 VSUBS xpredec0_bot_3v1024x8m81_0/nmos_5p04310591302066_3v1024x8m81_0/D
+ xpredec0_bot_3v1024x8m81_1/nmos_5p04310591302066_3v1024x8m81_0/D xpredec0_bot_3v1024x8m81_0/nmos_5p04310591302066_3v1024x8m81_0/D
+ A[0] vdd_uq2 xpredec0_bot_3v1024x8m81_1/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ xpredec0_bot_3v1024x8m81_0/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ xpredec0_bot_3v1024x8m81_0/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ nmos_5p04310591302040_3v1024x8m81_1/S pmos_5p04310591302069_3v1024x8m81_0/D vdd
+ vdd_uq2 VSUBS xpredec0_bot_3v1024x8m81
Xxpredec0_bot_3v1024x8m81_1 VSUBS xpredec0_bot_3v1024x8m81_1/nmos_5p04310591302066_3v1024x8m81_0/D
+ xpredec0_bot_3v1024x8m81_1/nmos_5p04310591302066_3v1024x8m81_0/D xpredec0_bot_3v1024x8m81_0/nmos_5p04310591302066_3v1024x8m81_0/D
+ A[1] vdd_uq2 xpredec0_bot_3v1024x8m81_1/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ xpredec0_bot_3v1024x8m81_0/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ xpredec0_bot_3v1024x8m81_1/pmos_1p2$$47504428_3v1024x8m81_0/pmos_5p04310591302063_3v1024x8m81_0/D
+ nmos_5p04310591302040_3v1024x8m81_1/S pmos_5p04310591302069_3v1024x8m81_0/D vdd
+ vdd_uq2 VSUBS xpredec0_bot_3v1024x8m81
X0 vdd_uq2 men a_3416_6773# vdd_uq2 pfet_03v3 ad=0.448p pd=2.72u as=0.162p ps=1.205u w=0.8u l=0.28u
X1 nmos_5p04310591302040_3v1024x8m81_1/S clk a_3091_6773# vdd_uq2 pfet_03v3 ad=0.218p pd=1.345u as=0.208p ps=1.32u w=0.8u l=0.28u
X2 a_3091_6773# men vdd_uq2 vdd_uq2 pfet_03v3 ad=0.208p pd=1.32u as=0.364p ps=2.51u w=0.8u l=0.28u
X3 a_3416_6773# clk nmos_5p04310591302040_3v1024x8m81_1/S vdd_uq2 pfet_03v3 ad=0.162p pd=1.205u as=0.218p ps=1.345u w=0.8u l=0.28u
.ends

.subckt prexdec_top_3v1024x8m81 A[6] A[4] xb[3] xc[2] xb[1] xb[2] xb[0] xa[1] xa[2]
+ xa[4] xa[5] xa[6] xa[7] A[0] A[3] A[5] A[1] xpredec1_3v1024x8m81_0/clk xpredec1_3v1024x8m81_0/pmos_1p2$$47109164_3v1024x8m81_0/pmos_5p04310591302062_3v1024x8m81_0/w_n202_n86#
+ xpredec1_3v1024x8m81_0/w_5024_6624# xa[0] A[2] xa[3] xc[1] xc[0] xpredec1_3v1024x8m81_0/xpredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/vdd
+ men xc[3] xpredec0_3v1024x8m81_1/vdd xpredec0_3v1024x8m81_1/clk VSUBS xpredec1_3v1024x8m81_0/vdd
Xxpredec1_3v1024x8m81_0 men xa[7] xa[6] xa[5] xa[4] xa[3] xa[2] xa[1] xa[0] xpredec1_3v1024x8m81_0/clk
+ xpredec1_3v1024x8m81_0/vdd xpredec1_3v1024x8m81_0/w_5024_6624# A[0] A[1] xpredec1_3v1024x8m81_0/vdd
+ xpredec0_3v1024x8m81_1/vdd A[2] VSUBS xpredec1_3v1024x8m81_0/xpredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/vdd
+ xpredec1_3v1024x8m81_0/pmos_1p2$$47109164_3v1024x8m81_0/pmos_5p04310591302062_3v1024x8m81_0/w_n202_n86#
+ xpredec1_3v1024x8m81
Xxpredec0_3v1024x8m81_0 xpredec0_3v1024x8m81_0/vss A[3] xb[1] xb[2] xb[3] A[4] xpredec0_3v1024x8m81_1/clk
+ xpredec0_3v1024x8m81_0/vss_uq0 xpredec0_3v1024x8m81_0/vdd_uq0 xpredec1_3v1024x8m81_0/vdd
+ xb[0] men xpredec0_3v1024x8m81_1/vdd VSUBS xpredec0_3v1024x8m81
Xxpredec0_3v1024x8m81_1 VSUBS A[5] xc[1] xc[2] xc[3] A[6] xpredec0_3v1024x8m81_1/clk
+ VSUBS xpredec0_3v1024x8m81_1/vdd xpredec1_3v1024x8m81_0/vdd xc[0] men xpredec0_3v1024x8m81_1/vdd
+ VSUBS xpredec0_3v1024x8m81
.ends

.subckt nmos_5p04310591302085_3v1024x8m81 D_uq1 D_uq0 a_530_n44# D a_n112_n44# a_209_n44#
+ a_369_n44# a_48_n44# S_uq1 S_uq0 S VSUBS
X0 D_uq1 a_n112_n44# S_uq1 VSUBS nfet_03v3 ad=1.2103p pd=5.175u as=2.0482p ps=10.19u w=4.655u l=0.28u
X1 S_uq0 a_369_n44# D VSUBS nfet_03v3 ad=1.22192p pd=5.18u as=1.2103p ps=5.175u w=4.655u l=0.28u
X2 D a_209_n44# S VSUBS nfet_03v3 ad=1.2103p pd=5.175u as=1.22192p ps=5.18u w=4.655u l=0.28u
X3 D_uq0 a_530_n44# S_uq0 VSUBS nfet_03v3 ad=2.0482p pd=10.19u as=1.22192p ps=5.18u w=4.655u l=0.28u
X4 S a_48_n44# D_uq1 VSUBS nfet_03v3 ad=1.22192p pd=5.18u as=1.2103p ps=5.175u w=4.655u l=0.28u
.ends

.subckt nmos_1p2$$48306220_3v1024x8m81 a_195_n34# a_355_n34# nmos_5p04310591302085_3v1024x8m81_0/S
+ a_n125_n34# nmos_5p04310591302085_3v1024x8m81_0/S_uq1 nmos_5p04310591302085_3v1024x8m81_0/S_uq0
+ a_34_n34# nmos_5p04310591302085_3v1024x8m81_0/D nmos_5p04310591302085_3v1024x8m81_0/D_uq1
+ nmos_5p04310591302085_3v1024x8m81_0/D_uq0 a_516_n34# VSUBS
Xnmos_5p04310591302085_3v1024x8m81_0 nmos_5p04310591302085_3v1024x8m81_0/D_uq1 nmos_5p04310591302085_3v1024x8m81_0/D_uq0
+ a_516_n34# nmos_5p04310591302085_3v1024x8m81_0/D a_n125_n34# a_195_n34# a_355_n34#
+ a_34_n34# nmos_5p04310591302085_3v1024x8m81_0/S_uq1 nmos_5p04310591302085_3v1024x8m81_0/S_uq0
+ nmos_5p04310591302085_3v1024x8m81_0/S VSUBS nmos_5p04310591302085_3v1024x8m81
.ends

.subckt pmos_5p04310591302092_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.1848p pd=1.72u as=0.1848p ps=1.72u w=0.42u l=0.465u
.ends

.subckt pmos_5p04310591302088_3v1024x8m81 D_uq2 D_uq1 D_uq0 D a_n252_n44# a_550_n44#
+ a_229_n44# w_n426_n86# S_uq4 S_uq2 S_uq3 S_uq1 a_390_n44# S_uq0 S a_n92_n44# a_1032_n44#
+ a_1192_n44# a_711_n44# a_69_n44# D_uq3 a_871_n44#
X0 D_uq1 a_390_n44# S_uq2 w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=1.52775p ps=6.345u w=5.82u l=0.28u
X1 D_uq3 a_n252_n44# S_uq4 w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=2.5608p ps=12.52u w=5.82u l=0.28u
X2 D_uq2 a_69_n44# S_uq3 w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=1.52775p ps=6.345u w=5.82u l=0.28u
X3 S_uq2 a_229_n44# D_uq2 w_n426_n86# pfet_03v3 ad=1.52775p pd=6.345u as=1.5132p ps=6.34u w=5.82u l=0.28u
X4 S_uq1 a_550_n44# D_uq1 w_n426_n86# pfet_03v3 ad=1.52775p pd=6.345u as=1.5132p ps=6.34u w=5.82u l=0.28u
X5 S_uq0 a_1192_n44# D_uq0 w_n426_n86# pfet_03v3 ad=2.5608p pd=12.52u as=1.5132p ps=6.34u w=5.82u l=0.28u
X6 D_uq0 a_1032_n44# S w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=1.52775p ps=6.345u w=5.82u l=0.28u
X7 S_uq3 a_n92_n44# D_uq3 w_n426_n86# pfet_03v3 ad=1.52775p pd=6.345u as=1.5132p ps=6.34u w=5.82u l=0.28u
X8 S a_871_n44# D w_n426_n86# pfet_03v3 ad=1.52775p pd=6.345u as=1.5132p ps=6.34u w=5.82u l=0.28u
X9 D a_711_n44# S_uq1 w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=1.52775p ps=6.345u w=5.82u l=0.28u
.ends

.subckt pmos_5p04310591302091_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=4.004p pd=19.08u as=4.004p ps=19.08u w=9.1u l=0.28u
.ends

.subckt pmos_1p2$$48624684_3v1024x8m81 pmos_5p04310591302091_3v1024x8m81_0/D a_n14_n34#
+ pmos_5p04310591302091_3v1024x8m81_0/S w_n133_n65#
Xpmos_5p04310591302091_3v1024x8m81_0 pmos_5p04310591302091_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302091_3v1024x8m81_0/S pmos_5p04310591302091_3v1024x8m81
.ends

.subckt pmos_1p2$$47330348_3v1024x8m81 pmos_5p04310591302041_3v1024x8m81_0/D a_n14_89#
+ pmos_5p04310591302041_3v1024x8m81_0/S w_n133_n65#
Xpmos_5p04310591302041_3v1024x8m81_0 pmos_5p04310591302041_3v1024x8m81_0/D a_n14_89#
+ w_n133_n65# pmos_5p04310591302041_3v1024x8m81_0/S pmos_5p04310591302041_3v1024x8m81
.ends

.subckt pmos_5p04310591302094_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.3872p pd=2.64u as=0.3872p ps=2.64u w=0.88u l=0.28u
.ends

.subckt nmos_5p04310591302093_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1576p pd=1.64u as=0.1576p ps=1.64u w=0.28u l=0.56u
.ends

.subckt nmos_5p04310591302090_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1576p pd=1.64u as=0.1576p ps=1.64u w=0.28u l=0.465u
.ends

.subckt pmos_5p04310591302087_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=4.6552p pd=22.04u as=4.6552p ps=22.04u w=10.58u l=0.28u
.ends

.subckt pmos_1p2$$47815724_3v1024x8m81 pmos_5p04310591302087_3v1024x8m81_0/S a_n14_n34#
+ pmos_5p04310591302087_3v1024x8m81_0/D w_n133_n65#
Xpmos_5p04310591302087_3v1024x8m81_0 pmos_5p04310591302087_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302087_3v1024x8m81_0/S pmos_5p04310591302087_3v1024x8m81
.ends

.subckt nmos_5p04310591302086_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.6182p pd=3.69u as=0.6182p ps=3.69u w=1.405u l=0.28u
.ends

.subckt nmos_1p2$$48302124_3v1024x8m81 nmos_5p04310591302086_3v1024x8m81_0/S nmos_5p04310591302086_3v1024x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p04310591302086_3v1024x8m81_0 nmos_5p04310591302086_3v1024x8m81_0/D a_n14_n34#
+ nmos_5p04310591302086_3v1024x8m81_0/S VSUBS nmos_5p04310591302086_3v1024x8m81
.ends

.subckt nmos_1p2$$48629804_3v1024x8m81 nmos_5p04310591302039_3v1024x8m81_0/S_uq0 nmos_5p04310591302039_3v1024x8m81_0/S
+ a_118_n34# nmos_5p04310591302039_3v1024x8m81_0/D a_n41_n34# VSUBS
Xnmos_5p04310591302039_3v1024x8m81_0 nmos_5p04310591302039_3v1024x8m81_0/D a_n41_n34#
+ a_118_n34# nmos_5p04310591302039_3v1024x8m81_0/S_uq0 nmos_5p04310591302039_3v1024x8m81_0/S
+ VSUBS nmos_5p04310591302039_3v1024x8m81
.ends

.subckt pmos_5p04310591302089_3v1024x8m81 D_uq2 D_uq1 a_2502_n44# D_uq0 a_1699_n44#
+ D a_n67_n44# a_2341_n44# a_1378_n44# a_2020_n44# a_1057_n44# a_n548_n44# S_uq9 S_uq8
+ S_uq7 S_uq6 a_94_n44# S_uq5 a_736_n44# a_n227_n44# S_uq4 S_uq2 S_uq3 a_896_n44#
+ S_uq1 S_uq0 w_n722_n86# S a_415_n44# a_2181_n44# a_1538_n44# a_575_n44# a_1860_n44#
+ D_uq8 D_uq7 a_1217_n44# a_n388_n44# D_uq6 a_254_n44# D_uq4 D_uq5 D_uq3
X0 D_uq8 a_n548_n44# S_uq9 w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=3.7708p ps=18.02u w=8.57u l=0.28u
X1 S_uq5 a_575_n44# D_uq5 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X2 D_uq5 a_415_n44# S_uq6 w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X3 D_uq3 a_1057_n44# S_uq4 w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X4 D a_2020_n44# S_uq1 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X5 S_uq4 a_896_n44# D_uq4 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X6 D_uq4 a_736_n44# S_uq5 w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X7 D_uq2 a_1378_n44# S_uq3 w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X8 D_uq0 a_2341_n44# S w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X9 S_uq7 a_n67_n44# D_uq7 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X10 D_uq1 a_1699_n44# S_uq2 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.24962p ps=9.095u w=8.57u l=0.28u
X11 S_uq0 a_2502_n44# D_uq0 w_n722_n86# pfet_03v3 ad=3.7708p pd=18.02u as=2.24962p ps=9.095u w=8.57u l=0.28u
X12 S_uq8 a_n388_n44# D_uq8 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X13 S_uq3 a_1217_n44# D_uq3 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X14 S_uq1 a_1860_n44# D_uq1 w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X15 S_uq2 a_1538_n44# D_uq2 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X16 S a_2181_n44# D w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X17 D_uq6 a_94_n44# S_uq7 w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X18 D_uq7 a_n227_n44# S_uq8 w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X19 S_uq6 a_254_n44# D_uq6 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
.ends

.subckt nmos_5p04310591302084_3v1024x8m81 D_uq2 D_uq1 D_uq0 a_1394_n44# D a_2357_n44#
+ a_1073_n44# a_2036_n44# a_n51_n44# a_1715_n44# a_752_n44# S_uq9 S_uq8 S_uq7 a_n532_n44#
+ S_uq6 S_uq5 a_431_n44# S_uq4 a_1554_n44# a_591_n44# S_uq2 S_uq3 a_2197_n44# S_uq1
+ a_n211_n44# S_uq0 S a_110_n44# a_1876_n44# a_1233_n44# a_270_n44# D_uq8 D_uq7 a_912_n44#
+ D_uq6 a_2518_n44# D_uq4 D_uq5 D_uq3 a_n372_n44# VSUBS
X0 S_uq6 a_270_n44# D_uq6 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X1 D_uq1 a_1715_n44# S_uq2 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.90167p ps=3.96u w=3.435u l=0.28u
X2 D_uq6 a_110_n44# S_uq7 VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X3 D a_2036_n44# S_uq1 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X4 S_uq7 a_n51_n44# D_uq7 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X5 S_uq5 a_591_n44# D_uq5 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X6 D_uq3 a_1073_n44# S_uq4 VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X7 D_uq5 a_431_n44# S_uq6 VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X8 D_uq0 a_2357_n44# S VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X9 D_uq2 a_1394_n44# S_uq3 VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X10 S_uq8 a_n372_n44# D_uq8 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X11 D_uq4 a_752_n44# S_uq5 VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X12 S_uq0 a_2518_n44# D_uq0 VSUBS nfet_03v3 ad=1.5114p pd=7.75u as=0.90167p ps=3.96u w=3.435u l=0.28u
X13 S_uq3 a_1233_n44# D_uq3 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X14 S_uq1 a_1876_n44# D_uq1 VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X15 D_uq7 a_n211_n44# S_uq8 VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X16 S a_2197_n44# D VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X17 S_uq2 a_1554_n44# D_uq2 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X18 D_uq8 a_n532_n44# S_uq9 VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=1.5114p ps=7.75u w=3.435u l=0.28u
X19 S_uq4 a_912_n44# D_uq4 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
.ends

.subckt nmos_1p2$$48308268_3v1024x8m81 nmos_5p04310591302084_3v1024x8m81_0/a_431_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/a_1073_n44# nmos_5p04310591302084_3v1024x8m81_0/a_591_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/a_2036_n44# nmos_5p04310591302084_3v1024x8m81_0/S_uq9
+ nmos_5p04310591302084_3v1024x8m81_0/a_110_n44# nmos_5p04310591302084_3v1024x8m81_0/a_1715_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/S_uq8 nmos_5p04310591302084_3v1024x8m81_0/a_270_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/S_uq7 nmos_5p04310591302084_3v1024x8m81_0/S_uq6
+ nmos_5p04310591302084_3v1024x8m81_0/a_n532_n44# nmos_5p04310591302084_3v1024x8m81_0/S_uq5
+ nmos_5p04310591302084_3v1024x8m81_0/S_uq4 nmos_5p04310591302084_3v1024x8m81_0/S_uq3
+ nmos_5p04310591302084_3v1024x8m81_0/a_912_n44# nmos_5p04310591302084_3v1024x8m81_0/a_1554_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/S_uq2 nmos_5p04310591302084_3v1024x8m81_0/S
+ nmos_5p04310591302084_3v1024x8m81_0/a_2197_n44# nmos_5p04310591302084_3v1024x8m81_0/S_uq1
+ nmos_5p04310591302084_3v1024x8m81_0/S_uq0 nmos_5p04310591302084_3v1024x8m81_0/a_n211_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/a_1233_n44# nmos_5p04310591302084_3v1024x8m81_0/a_1876_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/D_uq8 nmos_5p04310591302084_3v1024x8m81_0/D_uq7
+ nmos_5p04310591302084_3v1024x8m81_0/D_uq6 nmos_5p04310591302084_3v1024x8m81_0/D_uq5
+ nmos_5p04310591302084_3v1024x8m81_0/a_2518_n44# nmos_5p04310591302084_3v1024x8m81_0/D_uq4
+ nmos_5p04310591302084_3v1024x8m81_0/a_n51_n44# nmos_5p04310591302084_3v1024x8m81_0/D_uq3
+ nmos_5p04310591302084_3v1024x8m81_0/D_uq2 nmos_5p04310591302084_3v1024x8m81_0/a_n372_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/D_uq1 nmos_5p04310591302084_3v1024x8m81_0/D
+ nmos_5p04310591302084_3v1024x8m81_0/D_uq0 nmos_5p04310591302084_3v1024x8m81_0/a_752_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/a_1394_n44# nmos_5p04310591302084_3v1024x8m81_0/a_2357_n44#
+ VSUBS
Xnmos_5p04310591302084_3v1024x8m81_0 nmos_5p04310591302084_3v1024x8m81_0/D_uq2 nmos_5p04310591302084_3v1024x8m81_0/D_uq1
+ nmos_5p04310591302084_3v1024x8m81_0/D_uq0 nmos_5p04310591302084_3v1024x8m81_0/a_1394_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/D nmos_5p04310591302084_3v1024x8m81_0/a_2357_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/a_1073_n44# nmos_5p04310591302084_3v1024x8m81_0/a_2036_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/a_n51_n44# nmos_5p04310591302084_3v1024x8m81_0/a_1715_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/a_752_n44# nmos_5p04310591302084_3v1024x8m81_0/S_uq9
+ nmos_5p04310591302084_3v1024x8m81_0/S_uq8 nmos_5p04310591302084_3v1024x8m81_0/S_uq7
+ nmos_5p04310591302084_3v1024x8m81_0/a_n532_n44# nmos_5p04310591302084_3v1024x8m81_0/S_uq6
+ nmos_5p04310591302084_3v1024x8m81_0/S_uq5 nmos_5p04310591302084_3v1024x8m81_0/a_431_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/S_uq4 nmos_5p04310591302084_3v1024x8m81_0/a_1554_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/a_591_n44# nmos_5p04310591302084_3v1024x8m81_0/S_uq2
+ nmos_5p04310591302084_3v1024x8m81_0/S_uq3 nmos_5p04310591302084_3v1024x8m81_0/a_2197_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/S_uq1 nmos_5p04310591302084_3v1024x8m81_0/a_n211_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/S_uq0 nmos_5p04310591302084_3v1024x8m81_0/S
+ nmos_5p04310591302084_3v1024x8m81_0/a_110_n44# nmos_5p04310591302084_3v1024x8m81_0/a_1876_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/a_1233_n44# nmos_5p04310591302084_3v1024x8m81_0/a_270_n44#
+ nmos_5p04310591302084_3v1024x8m81_0/D_uq8 nmos_5p04310591302084_3v1024x8m81_0/D_uq7
+ nmos_5p04310591302084_3v1024x8m81_0/a_912_n44# nmos_5p04310591302084_3v1024x8m81_0/D_uq6
+ nmos_5p04310591302084_3v1024x8m81_0/a_2518_n44# nmos_5p04310591302084_3v1024x8m81_0/D_uq4
+ nmos_5p04310591302084_3v1024x8m81_0/D_uq5 nmos_5p04310591302084_3v1024x8m81_0/D_uq3
+ nmos_5p04310591302084_3v1024x8m81_0/a_n372_n44# VSUBS nmos_5p04310591302084_3v1024x8m81
.ends

.subckt nmos_5p04310591302083_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1646p pd=1.64u as=0.1646p ps=1.64u w=0.35u l=0.28u
.ends

.subckt pmos_5p04310591302074_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.1848p pd=1.72u as=0.1848p ps=1.72u w=0.42u l=0.56u
.ends

.subckt nmos_5p04310591302076_3v1024x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.28u
.ends

.subckt pmos_5p04310591302079_3v1024x8m81 D_uq2 D_uq1 D_uq0 D a_486_n44# a_165_n44#
+ a_n156_n44# S_uq2 S_uq1 S_uq0 S a_4_n44# a_646_n44# w_n330_n86# a_808_n44# a_325_n44#
X0 S_uq0 a_646_n44# D w_n330_n86# pfet_03v3 ad=0.27162p pd=1.555u as=0.2665p ps=1.545u w=1.025u l=0.28u
X1 D_uq1 a_165_n44# S_uq1 w_n330_n86# pfet_03v3 ad=0.2665p pd=1.545u as=0.26905p ps=1.55u w=1.025u l=0.28u
X2 D a_486_n44# S w_n330_n86# pfet_03v3 ad=0.2665p pd=1.545u as=0.26905p ps=1.55u w=1.025u l=0.28u
X3 S_uq1 a_4_n44# D_uq2 w_n330_n86# pfet_03v3 ad=0.26905p pd=1.55u as=0.2665p ps=1.545u w=1.025u l=0.28u
X4 D_uq2 a_n156_n44# S_uq2 w_n330_n86# pfet_03v3 ad=0.2665p pd=1.545u as=0.451p ps=2.93u w=1.025u l=0.28u
X5 S a_325_n44# D_uq1 w_n330_n86# pfet_03v3 ad=0.26905p pd=1.55u as=0.2665p ps=1.545u w=1.025u l=0.28u
X6 D_uq0 a_808_n44# S_uq0 w_n330_n86# pfet_03v3 ad=0.451p pd=2.93u as=0.27162p ps=1.555u w=1.025u l=0.28u
.ends

.subckt pmos_5p04310591302080_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.3445p pd=1.845u as=0.583p ps=3.53u w=1.325u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.583p pd=3.53u as=0.3445p ps=1.845u w=1.325u l=0.28u
.ends

.subckt nmos_5p04310591302078_3v1024x8m81 D_uq0 D S_uq0 S a_217_n44# a_n104_n44# a_56_n44#
+ VSUBS
X0 D_uq0 a_217_n44# S_uq0 VSUBS nfet_03v3 ad=0.4092p pd=2.74u as=0.24412p ps=1.455u w=0.93u l=0.28u
X1 S_uq0 a_56_n44# D VSUBS nfet_03v3 ad=0.24412p pd=1.455u as=0.2418p ps=1.45u w=0.93u l=0.28u
X2 D a_n104_n44# S VSUBS nfet_03v3 ad=0.2418p pd=1.45u as=0.4092p ps=2.74u w=0.93u l=0.28u
.ends

.subckt nmos_5p04310591302075_3v1024x8m81 D_uq2 D_uq1 D_uq0 D a_n252_n44# a_550_n44#
+ a_229_n44# S_uq4 S_uq2 S_uq3 S_uq1 a_390_n44# S_uq0 S a_n92_n44# a_1032_n44# a_1192_n44#
+ a_711_n44# a_69_n44# D_uq3 a_871_n44# VSUBS
X0 D_uq1 a_390_n44# S_uq2 VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.23492p ps=1.42u w=0.895u l=0.28u
X1 D_uq3 a_n252_n44# S_uq4 VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.3938p ps=2.67u w=0.895u l=0.28u
X2 D_uq2 a_69_n44# S_uq3 VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.23492p ps=1.42u w=0.895u l=0.28u
X3 S_uq2 a_229_n44# D_uq2 VSUBS nfet_03v3 ad=0.23492p pd=1.42u as=0.2327p ps=1.415u w=0.895u l=0.28u
X4 S_uq1 a_550_n44# D_uq1 VSUBS nfet_03v3 ad=0.23492p pd=1.42u as=0.2327p ps=1.415u w=0.895u l=0.28u
X5 S_uq0 a_1192_n44# D_uq0 VSUBS nfet_03v3 ad=0.3938p pd=2.67u as=0.2327p ps=1.415u w=0.895u l=0.28u
X6 D_uq0 a_1032_n44# S VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.23492p ps=1.42u w=0.895u l=0.28u
X7 S_uq3 a_n92_n44# D_uq3 VSUBS nfet_03v3 ad=0.23492p pd=1.42u as=0.2327p ps=1.415u w=0.895u l=0.28u
X8 S a_871_n44# D VSUBS nfet_03v3 ad=0.23492p pd=1.42u as=0.2327p ps=1.415u w=0.895u l=0.28u
X9 D a_711_n44# S_uq1 VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.23492p ps=1.42u w=0.895u l=0.28u
.ends

.subckt pmos_5p04310591302082_3v1024x8m81 a_20_n44# D_uq1 D_uq0 D a_181_n44# a_502_n44#
+ S_uq2 a_662_n44# S_uq1 a_n140_n44# S_uq0 S a_341_n44# w_n314_n86#
X0 S a_341_n44# D w_n314_n86# pfet_03v3 ad=0.30318p pd=1.68u as=0.3003p ps=1.675u w=1.155u l=0.28u
X1 S_uq0 a_662_n44# D_uq0 w_n314_n86# pfet_03v3 ad=0.5082p pd=3.19u as=0.3003p ps=1.675u w=1.155u l=0.28u
X2 D_uq0 a_502_n44# S w_n314_n86# pfet_03v3 ad=0.3003p pd=1.675u as=0.30318p ps=1.68u w=1.155u l=0.28u
X3 S_uq1 a_20_n44# D_uq1 w_n314_n86# pfet_03v3 ad=0.30318p pd=1.68u as=0.3003p ps=1.675u w=1.155u l=0.28u
X4 D a_181_n44# S_uq1 w_n314_n86# pfet_03v3 ad=0.3003p pd=1.675u as=0.30318p ps=1.68u w=1.155u l=0.28u
X5 D_uq1 a_n140_n44# S_uq2 w_n314_n86# pfet_03v3 ad=0.3003p pd=1.675u as=0.5082p ps=3.19u w=1.155u l=0.28u
.ends

.subckt nmos_5p04310591302081_3v1024x8m81 D_uq2 D_uq1 D_uq0 D a_634_n44# a_n168_n44#
+ a_313_n44# a_795_n44# S_uq2 a_474_n44# S_uq1 a_n8_n44# S_uq0 S a_153_n44# VSUBS
X0 D_uq1 a_153_n44# S_uq1 VSUBS nfet_03v3 ad=0.1079p pd=0.935u as=0.10892p ps=0.94u w=0.415u l=0.28u
X1 D a_474_n44# S VSUBS nfet_03v3 ad=0.1079p pd=0.935u as=0.10892p ps=0.94u w=0.415u l=0.28u
X2 D_uq2 a_n168_n44# S_uq2 VSUBS nfet_03v3 ad=0.1079p pd=0.935u as=0.1826p ps=1.71u w=0.415u l=0.28u
X3 S_uq1 a_n8_n44# D_uq2 VSUBS nfet_03v3 ad=0.10892p pd=0.94u as=0.1079p ps=0.935u w=0.415u l=0.28u
X4 D_uq0 a_795_n44# S_uq0 VSUBS nfet_03v3 ad=0.1826p pd=1.71u as=0.10892p ps=0.94u w=0.415u l=0.28u
X5 S a_313_n44# D_uq1 VSUBS nfet_03v3 ad=0.10892p pd=0.94u as=0.1079p ps=0.935u w=0.415u l=0.28u
X6 S_uq0 a_634_n44# D VSUBS nfet_03v3 ad=0.10892p pd=0.94u as=0.1079p ps=0.935u w=0.415u l=0.28u
.ends

.subckt pmos_5p04310591302077_3v1024x8m81 D_uq2 D_uq1 D_uq0 D a_n252_n44# a_550_n44#
+ a_229_n44# w_n426_n86# S_uq4 S_uq2 S_uq3 S_uq1 a_390_n44# S_uq0 S a_n92_n44# a_1032_n44#
+ a_1192_n44# a_711_n44# a_69_n44# D_uq3 a_871_n44#
X0 D_uq1 a_390_n44# S_uq2 w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.5775p ps=2.725u w=2.2u l=0.28u
X1 D_uq3 a_n252_n44# S_uq4 w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.968p ps=5.28u w=2.2u l=0.28u
X2 D_uq2 a_69_n44# S_uq3 w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.5775p ps=2.725u w=2.2u l=0.28u
X3 S_uq2 a_229_n44# D_uq2 w_n426_n86# pfet_03v3 ad=0.5775p pd=2.725u as=0.572p ps=2.72u w=2.2u l=0.28u
X4 S_uq1 a_550_n44# D_uq1 w_n426_n86# pfet_03v3 ad=0.5775p pd=2.725u as=0.572p ps=2.72u w=2.2u l=0.28u
X5 S_uq0 a_1192_n44# D_uq0 w_n426_n86# pfet_03v3 ad=0.968p pd=5.28u as=0.572p ps=2.72u w=2.2u l=0.28u
X6 D_uq0 a_1032_n44# S w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.5775p ps=2.725u w=2.2u l=0.28u
X7 S_uq3 a_n92_n44# D_uq3 w_n426_n86# pfet_03v3 ad=0.5775p pd=2.725u as=0.572p ps=2.72u w=2.2u l=0.28u
X8 S a_871_n44# D w_n426_n86# pfet_03v3 ad=0.5775p pd=2.725u as=0.572p ps=2.72u w=2.2u l=0.28u
X9 D a_711_n44# S_uq1 w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.5775p ps=2.725u w=2.2u l=0.28u
.ends

.subckt wen_v2_3v1024x8m81 IGWEN clk wen GWE vdd vss
Xnmos_5p04310591302076_3v1024x8m81_0 pmos_5p04310591302080_3v1024x8m81_0/D pmos_5p04310591302014_3v1024x8m81_2/S
+ pmos_5p04310591302014_3v1024x8m81_2/S vss vss vss nmos_5p04310591302076_3v1024x8m81
Xpmos_5p04310591302079_3v1024x8m81_0 pmos_5p04310591302079_3v1024x8m81_0/D pmos_5p04310591302079_3v1024x8m81_0/D
+ pmos_5p04310591302079_3v1024x8m81_0/D pmos_5p04310591302079_3v1024x8m81_0/D nmos_5p0431059130208_3v1024x8m81_1/S
+ nmos_5p0431059130208_3v1024x8m81_1/S nmos_5p0431059130208_3v1024x8m81_1/S vdd vdd
+ vdd vdd nmos_5p0431059130208_3v1024x8m81_1/S nmos_5p0431059130208_3v1024x8m81_1/S
+ vdd nmos_5p0431059130208_3v1024x8m81_1/S nmos_5p0431059130208_3v1024x8m81_1/S pmos_5p04310591302079_3v1024x8m81
Xpmos_5p04310591302080_3v1024x8m81_0 pmos_5p04310591302080_3v1024x8m81_0/D pmos_5p04310591302014_3v1024x8m81_2/S
+ pmos_5p04310591302014_3v1024x8m81_2/S vdd vdd vdd pmos_5p04310591302080_3v1024x8m81
Xnmos_5p0431059130208_3v1024x8m81_0 vss pmos_5p04310591302079_3v1024x8m81_0/D nmos_5p0431059130208_3v1024x8m81_1/D
+ vss nmos_5p0431059130208_3v1024x8m81
Xnmos_5p0431059130208_3v1024x8m81_1 nmos_5p0431059130208_3v1024x8m81_1/D nmos_5p0431059130208_3v1024x8m81_3/D
+ nmos_5p0431059130208_3v1024x8m81_1/S vss nmos_5p0431059130208_3v1024x8m81
Xnmos_1p2$$202595372_3v1024x8m81_0 pmos_5p04310591302014_3v1024x8m81_2/S vss pmos_5p04310591302041_3v1024x8m81_1/S
+ vss nmos_1p2$$202595372_3v1024x8m81
Xnmos_5p0431059130208_3v1024x8m81_2 vss wen nmos_5p0431059130208_3v1024x8m81_2/S vss
+ nmos_5p0431059130208_3v1024x8m81
Xnmos_1p2$$202595372_3v1024x8m81_1 pmos_5p04310591302041_3v1024x8m81_1/S pmos_5p04310591302041_3v1024x8m81_1/D
+ nmos_5p0431059130208_3v1024x8m81_4/D vss nmos_1p2$$202595372_3v1024x8m81
Xnmos_5p04310591302078_3v1024x8m81_0 pmos_5p04310591302082_3v1024x8m81_0/D pmos_5p04310591302082_3v1024x8m81_0/D
+ vss vss wen wen wen vss nmos_5p04310591302078_3v1024x8m81
Xnmos_5p0431059130208_3v1024x8m81_3 nmos_5p0431059130208_3v1024x8m81_3/D clk vss vss
+ nmos_5p0431059130208_3v1024x8m81
Xpmos_1p2$$202587180_3v1024x8m81_0 nmos_5p0431059130208_3v1024x8m81_4/D nmos_5p0431059130208_3v1024x8m81_2/S
+ pmos_5p04310591302041_3v1024x8m81_1/S vdd pmos_1p2$$202587180_3v1024x8m81
Xnmos_5p0431059130208_3v1024x8m81_4 nmos_5p0431059130208_3v1024x8m81_4/D nmos_5p0431059130208_3v1024x8m81_3/D
+ vss vss nmos_5p0431059130208_3v1024x8m81
Xnmos_5p04310591302075_3v1024x8m81_0 GWE GWE GWE GWE pmos_5p04310591302079_3v1024x8m81_0/D
+ pmos_5p04310591302079_3v1024x8m81_0/D pmos_5p04310591302079_3v1024x8m81_0/D vss
+ vss vss vss pmos_5p04310591302079_3v1024x8m81_0/D vss vss pmos_5p04310591302079_3v1024x8m81_0/D
+ pmos_5p04310591302079_3v1024x8m81_0/D pmos_5p04310591302079_3v1024x8m81_0/D pmos_5p04310591302079_3v1024x8m81_0/D
+ pmos_5p04310591302079_3v1024x8m81_0/D GWE pmos_5p04310591302079_3v1024x8m81_0/D
+ vss nmos_5p04310591302075_3v1024x8m81
Xnmos_5p04310591302075_3v1024x8m81_1 IGWEN IGWEN IGWEN IGWEN pmos_5p04310591302082_3v1024x8m81_0/D
+ pmos_5p04310591302082_3v1024x8m81_0/D pmos_5p04310591302082_3v1024x8m81_0/D vss
+ vss vss vss pmos_5p04310591302082_3v1024x8m81_0/D vss vss pmos_5p04310591302082_3v1024x8m81_0/D
+ pmos_5p04310591302082_3v1024x8m81_0/D pmos_5p04310591302082_3v1024x8m81_0/D pmos_5p04310591302082_3v1024x8m81_0/D
+ pmos_5p04310591302082_3v1024x8m81_0/D IGWEN pmos_5p04310591302082_3v1024x8m81_0/D
+ vss nmos_5p04310591302075_3v1024x8m81
Xpmos_5p04310591302082_3v1024x8m81_0 wen pmos_5p04310591302082_3v1024x8m81_0/D pmos_5p04310591302082_3v1024x8m81_0/D
+ pmos_5p04310591302082_3v1024x8m81_0/D wen wen vdd wen vdd wen vdd vdd wen vdd pmos_5p04310591302082_3v1024x8m81
Xpmos_1p2$$202586156_3v1024x8m81_0 pmos_5p04310591302014_3v1024x8m81_2/S pmos_5p04310591302041_3v1024x8m81_1/D
+ vdd vdd pmos_1p2$$202586156_3v1024x8m81
Xpmos_5p04310591302014_3v1024x8m81_0 vdd pmos_5p04310591302079_3v1024x8m81_0/D vdd
+ nmos_5p0431059130208_3v1024x8m81_1/D pmos_5p04310591302014_3v1024x8m81
Xpmos_5p04310591302014_3v1024x8m81_1 nmos_5p0431059130208_3v1024x8m81_3/D clk vdd
+ vdd pmos_5p04310591302014_3v1024x8m81
Xnmos_5p04310591302081_3v1024x8m81_0 pmos_5p04310591302079_3v1024x8m81_0/D pmos_5p04310591302079_3v1024x8m81_0/D
+ pmos_5p04310591302079_3v1024x8m81_0/D pmos_5p04310591302079_3v1024x8m81_0/D nmos_5p0431059130208_3v1024x8m81_1/S
+ nmos_5p0431059130208_3v1024x8m81_1/S nmos_5p0431059130208_3v1024x8m81_1/S nmos_5p0431059130208_3v1024x8m81_1/S
+ vss nmos_5p0431059130208_3v1024x8m81_1/S vss nmos_5p0431059130208_3v1024x8m81_1/S
+ vss vss nmos_5p0431059130208_3v1024x8m81_1/S vss nmos_5p04310591302081_3v1024x8m81
Xpmos_5p04310591302014_3v1024x8m81_2 vdd pmos_5p04310591302041_3v1024x8m81_1/S vdd
+ pmos_5p04310591302014_3v1024x8m81_2/S pmos_5p04310591302014_3v1024x8m81
Xnmos_1p2$$202596396_3v1024x8m81_0 pmos_5p04310591302041_3v1024x8m81_1/D vss pmos_5p04310591302014_3v1024x8m81_2/S
+ vss nmos_1p2$$202596396_3v1024x8m81
Xpmos_5p04310591302014_3v1024x8m81_3 vdd wen vdd nmos_5p0431059130208_3v1024x8m81_2/S
+ pmos_5p04310591302014_3v1024x8m81
Xpmos_5p04310591302014_3v1024x8m81_4 nmos_5p0431059130208_3v1024x8m81_4/D nmos_5p0431059130208_3v1024x8m81_3/D
+ vdd vdd pmos_5p04310591302014_3v1024x8m81
Xpmos_5p04310591302020_3v1024x8m81_0 pmos_5p04310591302080_3v1024x8m81_0/D nmos_5p0431059130208_3v1024x8m81_3/D
+ nmos_5p0431059130208_3v1024x8m81_3/D vdd nmos_5p0431059130208_3v1024x8m81_1/S nmos_5p0431059130208_3v1024x8m81_1/S
+ pmos_5p04310591302020_3v1024x8m81
Xnmos_5p04310591302010_3v1024x8m81_0 pmos_5p04310591302041_3v1024x8m81_1/S nmos_5p0431059130208_3v1024x8m81_3/D
+ nmos_5p0431059130208_3v1024x8m81_2/S vss nmos_5p04310591302010_3v1024x8m81
Xpmos_5p04310591302077_3v1024x8m81_0 IGWEN IGWEN IGWEN IGWEN pmos_5p04310591302082_3v1024x8m81_0/D
+ pmos_5p04310591302082_3v1024x8m81_0/D pmos_5p04310591302082_3v1024x8m81_0/D vdd
+ vdd vdd vdd vdd pmos_5p04310591302082_3v1024x8m81_0/D vdd vdd pmos_5p04310591302082_3v1024x8m81_0/D
+ pmos_5p04310591302082_3v1024x8m81_0/D pmos_5p04310591302082_3v1024x8m81_0/D pmos_5p04310591302082_3v1024x8m81_0/D
+ pmos_5p04310591302082_3v1024x8m81_0/D IGWEN pmos_5p04310591302082_3v1024x8m81_0/D
+ pmos_5p04310591302077_3v1024x8m81
Xpmos_5p04310591302041_3v1024x8m81_0 nmos_5p0431059130208_3v1024x8m81_1/D nmos_5p0431059130208_3v1024x8m81_4/D
+ vdd nmos_5p0431059130208_3v1024x8m81_1/S pmos_5p04310591302041_3v1024x8m81
Xpmos_5p04310591302041_3v1024x8m81_1 pmos_5p04310591302041_3v1024x8m81_1/D nmos_5p0431059130208_3v1024x8m81_3/D
+ vdd pmos_5p04310591302041_3v1024x8m81_1/S pmos_5p04310591302041_3v1024x8m81
Xpmos_5p04310591302077_3v1024x8m81_2 GWE GWE GWE GWE pmos_5p04310591302079_3v1024x8m81_0/D
+ pmos_5p04310591302079_3v1024x8m81_0/D pmos_5p04310591302079_3v1024x8m81_0/D vdd
+ vdd vdd vdd vdd pmos_5p04310591302079_3v1024x8m81_0/D vdd vdd pmos_5p04310591302079_3v1024x8m81_0/D
+ pmos_5p04310591302079_3v1024x8m81_0/D pmos_5p04310591302079_3v1024x8m81_0/D pmos_5p04310591302079_3v1024x8m81_0/D
+ pmos_5p04310591302079_3v1024x8m81_0/D GWE pmos_5p04310591302079_3v1024x8m81_0/D
+ pmos_5p04310591302077_3v1024x8m81
Xnmos_5p04310591302039_3v1024x8m81_0 pmos_5p04310591302080_3v1024x8m81_0/D nmos_5p0431059130208_3v1024x8m81_4/D
+ nmos_5p0431059130208_3v1024x8m81_4/D nmos_5p0431059130208_3v1024x8m81_1/S nmos_5p0431059130208_3v1024x8m81_1/S
+ vss nmos_5p04310591302039_3v1024x8m81
.ends

.subckt pmos_5p04310591302073_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.4563p pd=2.275u as=0.7722p ps=4.39u w=1.755u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.7722p pd=4.39u as=0.4563p ps=2.275u w=1.755u l=0.28u
.ends

.subckt pmos_1p2$$48623660_3v1024x8m81 a_n42_n34# w_n133_n66# pmos_5p04310591302073_3v1024x8m81_0/S
+ a_118_n34# pmos_5p04310591302073_3v1024x8m81_0/D pmos_5p04310591302073_3v1024x8m81_0/S_uq0
Xpmos_5p04310591302073_3v1024x8m81_0 pmos_5p04310591302073_3v1024x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302073_3v1024x8m81_0/S_uq0 pmos_5p04310591302073_3v1024x8m81_0/S
+ pmos_5p04310591302073_3v1024x8m81
.ends

.subckt gen_3v1024x8_3v1024x8m81 VSS tblhl cen clk WEN GWE wen_v2_3v1024x8m81_0/wen
+ VDD_uq3 VDD men pmos_5p04310591302088_3v1024x8m81_0/D IGWEN VDD_uq2
Xnmos_1p2$$48306220_3v1024x8m81_0 pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S
+ pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S VSS pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S
+ VSS VSS pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S pmos_5p04310591302088_3v1024x8m81_0/D
+ pmos_5p04310591302088_3v1024x8m81_0/D pmos_5p04310591302088_3v1024x8m81_0/D pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S
+ VSS nmos_1p2$$48306220_3v1024x8m81
Xnmos_1p2$$47342636_3v1024x8m81_0 nmos_1p2$$47342636_3v1024x8m81_1/nmos_5p04310591302053_3v1024x8m81_0/S
+ clk VSS VSS nmos_1p2$$47342636_3v1024x8m81
Xnmos_1p2$$47342636_3v1024x8m81_1 VSS men nmos_1p2$$47342636_3v1024x8m81_1/nmos_5p04310591302053_3v1024x8m81_0/S
+ VSS nmos_1p2$$47342636_3v1024x8m81
Xpmos_5p04310591302092_3v1024x8m81_0 pmos_5p04310591302092_3v1024x8m81_0/D pmos_5p04310591302074_3v1024x8m81_1/D
+ VDD VDD pmos_5p04310591302092_3v1024x8m81
Xpmos_5p04310591302088_3v1024x8m81_0 pmos_5p04310591302088_3v1024x8m81_0/D pmos_5p04310591302088_3v1024x8m81_0/D
+ pmos_5p04310591302088_3v1024x8m81_0/D pmos_5p04310591302088_3v1024x8m81_0/D pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S
+ pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S
+ VDD_uq3 VDD_uq3 VDD_uq3 VDD_uq3 VDD_uq3 pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S
+ VDD_uq3 VDD_uq3 pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S
+ pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S
+ pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S
+ pmos_5p04310591302088_3v1024x8m81_0/D pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S
+ pmos_5p04310591302088_3v1024x8m81
Xpmos_1p2$$48624684_3v1024x8m81_0 pmos_1p2$$48624684_3v1024x8m81_2/pmos_5p04310591302091_3v1024x8m81_0/S
+ pmos_5p04310591302051_3v1024x8m81_0/D VDD_uq2 VDD_uq2 pmos_1p2$$48624684_3v1024x8m81
Xpmos_1p2$$46273580_3v1024x8m81_0 VDD_uq2 pmos_5p04310591302051_3v1024x8m81_0/D VDD_uq2
+ pmos_5p04310591302051_3v1024x8m81_0/D pmos_1p2$$46273580_3v1024x8m81_0/pmos_5p0431059130203_3v1024x8m81_0/D
+ VDD_uq2 pmos_1p2$$46273580_3v1024x8m81
Xpmos_1p2$$48624684_3v1024x8m81_1 pmos_1p2$$48624684_3v1024x8m81_2/pmos_5p04310591302091_3v1024x8m81_0/S
+ pmos_1p2$$48623660_3v1024x8m81_0/pmos_5p04310591302073_3v1024x8m81_0/D VDD_uq2 VDD_uq2
+ pmos_1p2$$48624684_3v1024x8m81
Xpmos_1p2$$47330348_3v1024x8m81_0 pmos_1p2$$46273580_3v1024x8m81_0/pmos_5p0431059130203_3v1024x8m81_0/D
+ nmos_1p2$$47342636_3v1024x8m81_1/nmos_5p04310591302053_3v1024x8m81_0/S nmos_1p2$$46563372_3v1024x8m81_2/nmos_5p0431059130208_3v1024x8m81_0/S
+ VDD_uq2 pmos_1p2$$47330348_3v1024x8m81
Xpmos_5p04310591302094_3v1024x8m81_0 pmos_5p04310591302094_3v1024x8m81_0/D pmos_5p04310591302092_3v1024x8m81_0/D
+ VDD VDD pmos_5p04310591302094_3v1024x8m81
Xpmos_1p2$$48624684_3v1024x8m81_2 VDD_uq2 clk pmos_1p2$$48624684_3v1024x8m81_2/pmos_5p04310591302091_3v1024x8m81_0/S
+ VDD_uq2 pmos_1p2$$48624684_3v1024x8m81
Xnmos_5p04310591302093_3v1024x8m81_0 pmos_5p04310591302074_3v1024x8m81_0/D clk VSS
+ VSS nmos_5p04310591302093_3v1024x8m81
Xpmos_5p04310591302051_3v1024x8m81_0 pmos_5p04310591302051_3v1024x8m81_0/D nmos_1p2$$46563372_3v1024x8m81_2/nmos_5p0431059130208_3v1024x8m81_0/S
+ nmos_1p2$$46563372_3v1024x8m81_2/nmos_5p0431059130208_3v1024x8m81_0/S VDD_uq2 VDD_uq2
+ VDD_uq2 pmos_5p04310591302051_3v1024x8m81
Xnmos_5p04310591302093_3v1024x8m81_1 pmos_5p04310591302074_3v1024x8m81_1/D pmos_5p04310591302074_3v1024x8m81_0/D
+ VSS VSS nmos_5p04310591302093_3v1024x8m81
Xnmos_1p2$$46563372_3v1024x8m81_0 VSS nmos_1p2$$46563372_3v1024x8m81_0/nmos_5p0431059130208_3v1024x8m81_0/D
+ nmos_1p2$$47342636_3v1024x8m81_1/nmos_5p04310591302053_3v1024x8m81_0/S VSS nmos_1p2$$46563372_3v1024x8m81
Xnmos_1p2$$46563372_3v1024x8m81_1 pmos_1p2$$46273580_3v1024x8m81_0/pmos_5p0431059130203_3v1024x8m81_0/D
+ VSS pmos_5p04310591302051_3v1024x8m81_0/D VSS nmos_1p2$$46563372_3v1024x8m81
Xnmos_1p2$$46563372_3v1024x8m81_2 nmos_1p2$$46563372_3v1024x8m81_2/nmos_5p0431059130208_3v1024x8m81_0/S
+ pmos_1p2$$46273580_3v1024x8m81_0/pmos_5p0431059130203_3v1024x8m81_0/D nmos_1p2$$46563372_3v1024x8m81_0/nmos_5p0431059130208_3v1024x8m81_0/D
+ VSS nmos_1p2$$46563372_3v1024x8m81
Xnmos_5p04310591302090_3v1024x8m81_0 pmos_5p04310591302092_3v1024x8m81_0/D pmos_5p04310591302074_3v1024x8m81_1/D
+ VSS VSS nmos_5p04310591302090_3v1024x8m81
Xpmos_1p2$$47815724_3v1024x8m81_0 pmos_1p2$$47815724_3v1024x8m81_3/pmos_5p04310591302087_3v1024x8m81_0/S
+ tblhl VDD_uq2 VDD_uq2 pmos_1p2$$47815724_3v1024x8m81
Xpmos_1p2$$46285868_3v1024x8m81_0 VDD_uq2 VDD_uq2 nmos_1p2$$47342636_3v1024x8m81_1/nmos_5p04310591302053_3v1024x8m81_0/S
+ nmos_1p2$$46563372_3v1024x8m81_0/nmos_5p0431059130208_3v1024x8m81_0/D pmos_1p2$$46285868_3v1024x8m81
Xpmos_1p2$$46285868_3v1024x8m81_1 VDD_uq2 nmos_1p2$$46563372_3v1024x8m81_2/nmos_5p0431059130208_3v1024x8m81_0/S
+ nmos_1p2$$46563372_3v1024x8m81_0/nmos_5p0431059130208_3v1024x8m81_0/D cen pmos_1p2$$46285868_3v1024x8m81
Xpmos_1p2$$47815724_3v1024x8m81_1 VDD_uq2 pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S
+ pmos_1p2$$47815724_3v1024x8m81_3/pmos_5p04310591302087_3v1024x8m81_0/S VDD_uq2 pmos_1p2$$47815724_3v1024x8m81
Xpmos_1p2$$47815724_3v1024x8m81_2 VDD_uq2 tblhl pmos_1p2$$47815724_3v1024x8m81_3/pmos_5p04310591302087_3v1024x8m81_0/S
+ VDD_uq2 pmos_1p2$$47815724_3v1024x8m81
Xnmos_1p2$$48302124_3v1024x8m81_0 VSS pmos_1p2$$48623660_3v1024x8m81_0/pmos_5p04310591302073_3v1024x8m81_0/D
+ pmos_5p04310591302094_3v1024x8m81_0/D VSS nmos_1p2$$48302124_3v1024x8m81
Xpmos_1p2$$47815724_3v1024x8m81_3 pmos_1p2$$47815724_3v1024x8m81_3/pmos_5p04310591302087_3v1024x8m81_0/S
+ pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S VDD_uq2 VDD_uq2
+ pmos_1p2$$47815724_3v1024x8m81
Xnmos_1p2$$48629804_3v1024x8m81_0 VSS VSS nmos_1p2$$46563372_3v1024x8m81_2/nmos_5p0431059130208_3v1024x8m81_0/S
+ pmos_5p04310591302051_3v1024x8m81_0/D nmos_1p2$$46563372_3v1024x8m81_2/nmos_5p0431059130208_3v1024x8m81_0/S
+ VSS nmos_1p2$$48629804_3v1024x8m81
Xpmos_1p2$$47815724_3v1024x8m81_4 VDD_uq2 pmos_1p2$$47815724_3v1024x8m81_3/pmos_5p04310591302087_3v1024x8m81_0/S
+ pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S VDD_uq2 pmos_1p2$$47815724_3v1024x8m81
Xpmos_5p04310591302089_3v1024x8m81_0 men men pmos_5p04310591302088_3v1024x8m81_0/D
+ men pmos_5p04310591302088_3v1024x8m81_0/D men pmos_5p04310591302088_3v1024x8m81_0/D
+ pmos_5p04310591302088_3v1024x8m81_0/D pmos_5p04310591302088_3v1024x8m81_0/D pmos_5p04310591302088_3v1024x8m81_0/D
+ pmos_5p04310591302088_3v1024x8m81_0/D pmos_5p04310591302088_3v1024x8m81_0/D VDD_uq3
+ VDD_uq3 VDD_uq3 VDD_uq3 pmos_5p04310591302088_3v1024x8m81_0/D VDD_uq3 pmos_5p04310591302088_3v1024x8m81_0/D
+ pmos_5p04310591302088_3v1024x8m81_0/D VDD_uq3 VDD_uq3 VDD_uq3 pmos_5p04310591302088_3v1024x8m81_0/D
+ VDD_uq3 VDD_uq3 VDD_uq3 VDD_uq3 pmos_5p04310591302088_3v1024x8m81_0/D pmos_5p04310591302088_3v1024x8m81_0/D
+ pmos_5p04310591302088_3v1024x8m81_0/D pmos_5p04310591302088_3v1024x8m81_0/D pmos_5p04310591302088_3v1024x8m81_0/D
+ men men pmos_5p04310591302088_3v1024x8m81_0/D pmos_5p04310591302088_3v1024x8m81_0/D
+ men pmos_5p04310591302088_3v1024x8m81_0/D men men men pmos_5p04310591302089_3v1024x8m81
Xnmos_1p2$$48308268_3v1024x8m81_0 pmos_5p04310591302088_3v1024x8m81_0/D pmos_5p04310591302088_3v1024x8m81_0/D
+ pmos_5p04310591302088_3v1024x8m81_0/D pmos_5p04310591302088_3v1024x8m81_0/D VSS
+ pmos_5p04310591302088_3v1024x8m81_0/D pmos_5p04310591302088_3v1024x8m81_0/D VSS
+ pmos_5p04310591302088_3v1024x8m81_0/D VSS VSS pmos_5p04310591302088_3v1024x8m81_0/D
+ VSS VSS VSS pmos_5p04310591302088_3v1024x8m81_0/D pmos_5p04310591302088_3v1024x8m81_0/D
+ VSS VSS pmos_5p04310591302088_3v1024x8m81_0/D VSS VSS pmos_5p04310591302088_3v1024x8m81_0/D
+ pmos_5p04310591302088_3v1024x8m81_0/D pmos_5p04310591302088_3v1024x8m81_0/D men
+ men men men pmos_5p04310591302088_3v1024x8m81_0/D men pmos_5p04310591302088_3v1024x8m81_0/D
+ men men pmos_5p04310591302088_3v1024x8m81_0/D men men men pmos_5p04310591302088_3v1024x8m81_0/D
+ pmos_5p04310591302088_3v1024x8m81_0/D pmos_5p04310591302088_3v1024x8m81_0/D VSS
+ nmos_1p2$$48308268_3v1024x8m81
Xpmos_1p2$$47815724_3v1024x8m81_5 VDD_uq2 pmos_1p2$$48624684_3v1024x8m81_2/pmos_5p04310591302091_3v1024x8m81_0/S
+ pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S VDD_uq2 pmos_1p2$$47815724_3v1024x8m81
Xnmos_5p04310591302083_3v1024x8m81_0 pmos_5p04310591302094_3v1024x8m81_0/D pmos_5p04310591302092_3v1024x8m81_0/D
+ VSS VSS nmos_5p04310591302083_3v1024x8m81
Xnmos_1p2$$46551084_3v1024x8m81_0 cen nmos_1p2$$47342636_3v1024x8m81_1/nmos_5p04310591302053_3v1024x8m81_0/S
+ nmos_1p2$$46563372_3v1024x8m81_2/nmos_5p0431059130208_3v1024x8m81_0/S VSS nmos_1p2$$46551084_3v1024x8m81
Xpmos_1p2$$47815724_3v1024x8m81_6 pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S
+ pmos_1p2$$47815724_3v1024x8m81_3/pmos_5p04310591302087_3v1024x8m81_0/S VDD_uq2 VDD_uq2
+ pmos_1p2$$47815724_3v1024x8m81
Xpmos_1p2$$47815724_3v1024x8m81_7 pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S
+ pmos_1p2$$48624684_3v1024x8m81_2/pmos_5p04310591302091_3v1024x8m81_0/S VDD_uq2 VDD_uq2
+ pmos_1p2$$47815724_3v1024x8m81
Xpmos_5p04310591302074_3v1024x8m81_0 pmos_5p04310591302074_3v1024x8m81_0/D clk VDD
+ VDD pmos_5p04310591302074_3v1024x8m81
Xwen_v2_3v1024x8m81_0 IGWEN clk wen_v2_3v1024x8m81_0/wen GWE VDD VSS wen_v2_3v1024x8m81
Xpmos_5p04310591302074_3v1024x8m81_1 pmos_5p04310591302074_3v1024x8m81_1/D pmos_5p04310591302074_3v1024x8m81_0/D
+ VDD VDD pmos_5p04310591302074_3v1024x8m81
Xpmos_1p2$$48623660_3v1024x8m81_0 pmos_5p04310591302094_3v1024x8m81_0/D VDD VDD pmos_5p04310591302094_3v1024x8m81_0/D
+ pmos_1p2$$48623660_3v1024x8m81_0/pmos_5p04310591302073_3v1024x8m81_0/D VDD pmos_1p2$$48623660_3v1024x8m81
X0 a_8790_2243# tblhl pmos_1p2$$47815724_3v1024x8m81_3/pmos_5p04310591302087_3v1024x8m81_0/S VSS nfet_03v3 ad=0.5499p pd=2.635u as=0.5499p ps=2.635u w=2.115u l=0.28u
X1 a_3606_4291# men VDD_uq2 VDD_uq2 pfet_03v3 ad=0.2769p pd=1.585u as=0.50587p ps=3.08u w=1.065u l=0.28u
X2 a_7891_338# pmos_1p2$$48624684_3v1024x8m81_2/pmos_5p04310591302091_3v1024x8m81_0/S pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S VSS nfet_03v3 ad=2.2009p pd=8.985u as=2.2009p ps=8.985u w=8.465u l=0.28u
X3 a_6888_183# clk a_6728_183# VSS nfet_03v3 ad=2.7521p pd=11.105u as=2.7521p ps=11.105u w=10.585u l=0.28u
X4 VSS pmos_1p2$$47815724_3v1024x8m81_3/pmos_5p04310591302087_3v1024x8m81_0/S a_7891_338# VSS nfet_03v3 ad=3.93622p pd=17.86u as=2.2009p ps=8.985u w=8.465u l=0.28u
X5 pmos_1p2$$47815724_3v1024x8m81_3/pmos_5p04310591302087_3v1024x8m81_0/S tblhl a_8470_2243# VSS nfet_03v3 ad=0.5499p pd=2.635u as=0.5499p ps=2.635u w=2.115u l=0.28u
X6 a_8470_2243# pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S VSS VSS nfet_03v3 ad=0.5499p pd=2.635u as=0.96232p ps=5.14u w=2.115u l=0.28u
X7 pmos_1p2$$48624684_3v1024x8m81_2/pmos_5p04310591302091_3v1024x8m81_0/S pmos_5p04310591302051_3v1024x8m81_0/D a_6888_183# VSS nfet_03v3 ad=5.2925p pd=22.17u as=2.7521p ps=11.105u w=10.585u l=0.28u
X8 a_7571_338# pmos_1p2$$47815724_3v1024x8m81_3/pmos_5p04310591302087_3v1024x8m81_0/S VSS VSS nfet_03v3 ad=2.2009p pd=8.985u as=3.85157p ps=17.84u w=8.465u l=0.28u
X9 pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S pmos_1p2$$48624684_3v1024x8m81_2/pmos_5p04310591302091_3v1024x8m81_0/S a_7571_338# VSS nfet_03v3 ad=2.2009p pd=8.985u as=2.2009p ps=8.985u w=8.465u l=0.28u
X10 a_6728_183# pmos_1p2$$48623660_3v1024x8m81_0/pmos_5p04310591302073_3v1024x8m81_0/D VSS VSS nfet_03v3 ad=2.7521p pd=11.105u as=4.6574p ps=22.05u w=10.585u l=0.28u
X11 nmos_1p2$$47342636_3v1024x8m81_1/nmos_5p04310591302053_3v1024x8m81_0/S clk a_3606_4291# VDD_uq2 pfet_03v3 ad=0.50587p pd=3.08u as=0.2769p ps=1.585u w=1.065u l=0.28u
X12 VSS pmos_1p2$$47815724_3v1024x8m81_7/pmos_5p04310591302087_3v1024x8m81_0/S a_8790_2243# VSS nfet_03v3 ad=0.99405p pd=5.17u as=0.5499p ps=2.635u w=2.115u l=0.28u
.ends

.subckt pmos_5p04310591302055_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=4.1052p pd=19.54u as=4.1052p ps=19.54u w=9.33u l=0.28u
.ends

.subckt nmos_5p04310591302054_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.8634p pd=9.35u as=1.8634p ps=9.35u w=4.235u l=0.28u
.ends

.subckt ypredec1_ys_3v1024x8m81 pmos_5p04310591302055_3v1024x8m81_1/S a_187_1127#
+ pmos_5p04310591302055_3v1024x8m81_3/S nmos_5p04310591302054_3v1024x8m81_3/D pmos_5p04310591302055_3v1024x8m81_3/D
+ VSUBS
Xpmos_5p04310591302055_3v1024x8m81_0 pmos_5p04310591302055_3v1024x8m81_0/D a_187_1127#
+ pmos_5p04310591302055_3v1024x8m81_3/D pmos_5p04310591302055_3v1024x8m81_3/D pmos_5p04310591302055_3v1024x8m81
Xpmos_5p04310591302055_3v1024x8m81_1 pmos_5p04310591302055_3v1024x8m81_3/D pmos_5p04310591302055_3v1024x8m81_0/D
+ pmos_5p04310591302055_3v1024x8m81_3/D pmos_5p04310591302055_3v1024x8m81_1/S pmos_5p04310591302055_3v1024x8m81
Xpmos_5p04310591302055_3v1024x8m81_2 pmos_5p04310591302055_3v1024x8m81_3/S pmos_5p04310591302055_3v1024x8m81_0/D
+ pmos_5p04310591302055_3v1024x8m81_3/D pmos_5p04310591302055_3v1024x8m81_3/D pmos_5p04310591302055_3v1024x8m81
Xpmos_5p04310591302055_3v1024x8m81_3 pmos_5p04310591302055_3v1024x8m81_3/D pmos_5p04310591302055_3v1024x8m81_0/D
+ pmos_5p04310591302055_3v1024x8m81_3/D pmos_5p04310591302055_3v1024x8m81_3/S pmos_5p04310591302055_3v1024x8m81
Xnmos_5p04310591302054_3v1024x8m81_0 pmos_5p04310591302055_3v1024x8m81_3/S pmos_5p04310591302055_3v1024x8m81_0/D
+ nmos_5p04310591302054_3v1024x8m81_3/D VSUBS nmos_5p04310591302054_3v1024x8m81
Xnmos_5p04310591302054_3v1024x8m81_1 nmos_5p04310591302054_3v1024x8m81_3/D pmos_5p04310591302055_3v1024x8m81_0/D
+ pmos_5p04310591302055_3v1024x8m81_1/S VSUBS nmos_5p04310591302054_3v1024x8m81
Xnmos_5p04310591302054_3v1024x8m81_2 pmos_5p04310591302055_3v1024x8m81_0/D a_187_1127#
+ nmos_5p04310591302054_3v1024x8m81_3/D VSUBS nmos_5p04310591302054_3v1024x8m81
Xnmos_5p04310591302054_3v1024x8m81_3 nmos_5p04310591302054_3v1024x8m81_3/D pmos_5p04310591302055_3v1024x8m81_0/D
+ pmos_5p04310591302055_3v1024x8m81_3/S VSUBS nmos_5p04310591302054_3v1024x8m81
.ends

.subckt pmos_5p04310591302060_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=1.1638p pd=6.17u as=1.1638p ps=6.17u w=2.645u l=0.28u
.ends

.subckt pmos_1p2$$47821868_3v1024x8m81 pmos_5p04310591302060_3v1024x8m81_0/S w_n133_n66#
+ a_n14_n34# pmos_5p04310591302060_3v1024x8m81_0/D
Xpmos_5p04310591302060_3v1024x8m81_0 pmos_5p04310591302060_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302060_3v1024x8m81_0/S pmos_5p04310591302060_3v1024x8m81
.ends

.subckt pmos_5p04310591302061_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=1.1836p pd=6.26u as=1.1836p ps=6.26u w=2.69u l=0.28u
.ends

.subckt pmos_1p2$$47820844_3v1024x8m81 pmos_5p04310591302061_3v1024x8m81_0/S a_n14_n34#
+ pmos_5p04310591302061_3v1024x8m81_0/D w_n133_n65#
Xpmos_5p04310591302061_3v1024x8m81_0 pmos_5p04310591302061_3v1024x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302061_3v1024x8m81_0/S pmos_5p04310591302061_3v1024x8m81
.ends

.subckt ypredec1_xa_3v1024x8m81 m1_n40_n2861# pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ a_145_n4683# m3_0_n4986# pmos_1p2$$47820844_3v1024x8m81_2/w_n133_n65# M3_M2$$47819820_3v1024x8m81_0/VSUBS
+ m1_n40_n3567# m1_n40_n3285# a_0_56# a_465_n4683# m1_n40_n3426# m1_n40_n3144# m1_n40_n3003#
+ a_305_n4683# pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/S
+ pmos_1p2$$47821868_3v1024x8m81_3/w_n133_n66#
Xpmos_1p2$$47821868_3v1024x8m81_0 pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/S
+ pmos_1p2$$47821868_3v1024x8m81_3/w_n133_n66# a_145_n4683# pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/D
+ pmos_1p2$$47821868_3v1024x8m81
Xpmos_1p2$$47821868_3v1024x8m81_2 pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/D
+ pmos_1p2$$47821868_3v1024x8m81_3/w_n133_n66# a_305_n4683# pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/S
+ pmos_1p2$$47821868_3v1024x8m81
Xpmos_1p2$$47821868_3v1024x8m81_3 pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/S
+ pmos_1p2$$47821868_3v1024x8m81_3/w_n133_n66# a_465_n4683# pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/D
+ pmos_1p2$$47821868_3v1024x8m81
Xpmos_1p2$$47820844_3v1024x8m81_0 pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/S
+ pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/D pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ pmos_1p2$$47820844_3v1024x8m81_2/w_n133_n65# pmos_1p2$$47820844_3v1024x8m81
Xpmos_1p2$$47820844_3v1024x8m81_1 pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/D pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/S
+ pmos_1p2$$47820844_3v1024x8m81_2/w_n133_n65# pmos_1p2$$47820844_3v1024x8m81
Xpmos_1p2$$47820844_3v1024x8m81_2 pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/S
+ pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/D pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ pmos_1p2$$47820844_3v1024x8m81_2/w_n133_n65# pmos_1p2$$47820844_3v1024x8m81
Xnmos_1p2$$46551084_3v1024x8m81_0 M3_M2$$47819820_3v1024x8m81_0/VSUBS pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/D
+ pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D M3_M2$$47819820_3v1024x8m81_0/VSUBS
+ nmos_1p2$$46551084_3v1024x8m81
Xnmos_1p2$$46551084_3v1024x8m81_1 pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/D M3_M2$$47819820_3v1024x8m81_0/VSUBS
+ M3_M2$$47819820_3v1024x8m81_0/VSUBS nmos_1p2$$46551084_3v1024x8m81
Xnmos_1p2$$46551084_3v1024x8m81_2 pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/D M3_M2$$47819820_3v1024x8m81_0/VSUBS
+ M3_M2$$47819820_3v1024x8m81_0/VSUBS nmos_1p2$$46551084_3v1024x8m81
X0 a_361_n4624# a_305_n4683# a_201_n4624# M3_M2$$47819820_3v1024x8m81_0/VSUBS nfet_03v3 ad=0.8268p pd=3.7u as=0.8268p ps=3.7u w=3.18u l=0.28u
X1 a_201_n4624# a_145_n4683# M3_M2$$47819820_3v1024x8m81_0/VSUBS M3_M2$$47819820_3v1024x8m81_0/VSUBS nfet_03v3 ad=0.8268p pd=3.7u as=1.4469p ps=7.27u w=3.18u l=0.28u
X2 pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/D a_465_n4683# a_361_n4624# M3_M2$$47819820_3v1024x8m81_0/VSUBS nfet_03v3 ad=1.5423p pd=7.33u as=0.8268p ps=3.7u w=3.18u l=0.28u
.ends

.subckt ypredec1_xax8_3v1024x8m81 ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xa_3v1024x8m81_6/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xa_3v1024x8m81_5/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xa_3v1024x8m81_3/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xa_3v1024x8m81_4/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xa_3v1024x8m81_5/a_0_56# ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/w_n133_n66#
+ ypredec1_xa_3v1024x8m81_0/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xa_3v1024x8m81_1/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xa_3v1024x8m81_2/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xa_3v1024x8m81_7/a_145_n4683# ypredec1_xa_3v1024x8m81_5/a_465_n4683# ypredec1_xa_3v1024x8m81_6/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_3/a_145_n4683# ypredec1_xa_3v1024x8m81_7/a_305_n4683# ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/S
+ ypredec1_xa_3v1024x8m81_7/a_465_n4683# ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47820844_3v1024x8m81_2/w_n133_n65#
+ VSUBS
Xypredec1_xa_3v1024x8m81_0 ypredec1_xa_3v1024x8m81_7/a_465_n4683# ypredec1_xa_3v1024x8m81_0/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xa_3v1024x8m81_3/a_145_n4683# VSUBS ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47820844_3v1024x8m81_2/w_n133_n65#
+ VSUBS ypredec1_xa_3v1024x8m81_7/a_145_n4683# ypredec1_xa_3v1024x8m81_5/a_465_n4683#
+ ypredec1_xa_3v1024x8m81_0/a_0_56# ypredec1_xa_3v1024x8m81_5/a_465_n4683# ypredec1_xa_3v1024x8m81_6/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_3/a_145_n4683# ypredec1_xa_3v1024x8m81_7/a_305_n4683# ypredec1_xa_3v1024x8m81_7/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/S
+ ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/w_n133_n66# ypredec1_xa_3v1024x8m81
Xypredec1_xa_3v1024x8m81_1 ypredec1_xa_3v1024x8m81_7/a_465_n4683# ypredec1_xa_3v1024x8m81_1/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xa_3v1024x8m81_3/a_145_n4683# VSUBS ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47820844_3v1024x8m81_2/w_n133_n65#
+ VSUBS ypredec1_xa_3v1024x8m81_7/a_145_n4683# ypredec1_xa_3v1024x8m81_5/a_465_n4683#
+ ypredec1_xa_3v1024x8m81_5/a_0_56# ypredec1_xa_3v1024x8m81_5/a_465_n4683# ypredec1_xa_3v1024x8m81_6/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_3/a_145_n4683# ypredec1_xa_3v1024x8m81_7/a_305_n4683# ypredec1_xa_3v1024x8m81_6/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/S
+ ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/w_n133_n66# ypredec1_xa_3v1024x8m81
Xypredec1_xa_3v1024x8m81_2 ypredec1_xa_3v1024x8m81_7/a_465_n4683# ypredec1_xa_3v1024x8m81_2/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xa_3v1024x8m81_3/a_145_n4683# VSUBS ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47820844_3v1024x8m81_2/w_n133_n65#
+ VSUBS ypredec1_xa_3v1024x8m81_7/a_145_n4683# ypredec1_xa_3v1024x8m81_5/a_465_n4683#
+ VSUBS ypredec1_xa_3v1024x8m81_7/a_465_n4683# ypredec1_xa_3v1024x8m81_6/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_3/a_145_n4683# ypredec1_xa_3v1024x8m81_7/a_305_n4683# ypredec1_xa_3v1024x8m81_6/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/S
+ ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/w_n133_n66# ypredec1_xa_3v1024x8m81
Xypredec1_xa_3v1024x8m81_3 ypredec1_xa_3v1024x8m81_7/a_465_n4683# ypredec1_xa_3v1024x8m81_3/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xa_3v1024x8m81_3/a_145_n4683# VSUBS ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47820844_3v1024x8m81_2/w_n133_n65#
+ VSUBS ypredec1_xa_3v1024x8m81_7/a_145_n4683# ypredec1_xa_3v1024x8m81_5/a_465_n4683#
+ ypredec1_xa_3v1024x8m81_3/a_0_56# ypredec1_xa_3v1024x8m81_7/a_465_n4683# ypredec1_xa_3v1024x8m81_6/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_3/a_145_n4683# ypredec1_xa_3v1024x8m81_7/a_305_n4683# ypredec1_xa_3v1024x8m81_7/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/S
+ ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/w_n133_n66# ypredec1_xa_3v1024x8m81
Xypredec1_xa_3v1024x8m81_4 ypredec1_xa_3v1024x8m81_7/a_465_n4683# ypredec1_xa_3v1024x8m81_4/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xa_3v1024x8m81_7/a_145_n4683# VSUBS ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47820844_3v1024x8m81_2/w_n133_n65#
+ VSUBS ypredec1_xa_3v1024x8m81_7/a_145_n4683# ypredec1_xa_3v1024x8m81_5/a_465_n4683#
+ ypredec1_xa_3v1024x8m81_4/a_0_56# ypredec1_xa_3v1024x8m81_5/a_465_n4683# ypredec1_xa_3v1024x8m81_6/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_3/a_145_n4683# ypredec1_xa_3v1024x8m81_7/a_305_n4683# ypredec1_xa_3v1024x8m81_7/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/S
+ ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/w_n133_n66# ypredec1_xa_3v1024x8m81
Xypredec1_xa_3v1024x8m81_5 ypredec1_xa_3v1024x8m81_7/a_465_n4683# ypredec1_xa_3v1024x8m81_5/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xa_3v1024x8m81_7/a_145_n4683# VSUBS ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47820844_3v1024x8m81_2/w_n133_n65#
+ VSUBS ypredec1_xa_3v1024x8m81_7/a_145_n4683# ypredec1_xa_3v1024x8m81_5/a_465_n4683#
+ ypredec1_xa_3v1024x8m81_5/a_0_56# ypredec1_xa_3v1024x8m81_5/a_465_n4683# ypredec1_xa_3v1024x8m81_6/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_3/a_145_n4683# ypredec1_xa_3v1024x8m81_7/a_305_n4683# ypredec1_xa_3v1024x8m81_6/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/S
+ ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/w_n133_n66# ypredec1_xa_3v1024x8m81
Xypredec1_xa_3v1024x8m81_6 ypredec1_xa_3v1024x8m81_7/a_465_n4683# ypredec1_xa_3v1024x8m81_6/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xa_3v1024x8m81_7/a_145_n4683# VSUBS ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47820844_3v1024x8m81_2/w_n133_n65#
+ VSUBS ypredec1_xa_3v1024x8m81_7/a_145_n4683# ypredec1_xa_3v1024x8m81_5/a_465_n4683#
+ ypredec1_xa_3v1024x8m81_6/a_0_56# ypredec1_xa_3v1024x8m81_7/a_465_n4683# ypredec1_xa_3v1024x8m81_6/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_3/a_145_n4683# ypredec1_xa_3v1024x8m81_7/a_305_n4683# ypredec1_xa_3v1024x8m81_6/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/S
+ ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/w_n133_n66# ypredec1_xa_3v1024x8m81
Xypredec1_xa_3v1024x8m81_7 ypredec1_xa_3v1024x8m81_7/a_465_n4683# ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xa_3v1024x8m81_7/a_145_n4683# VSUBS ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47820844_3v1024x8m81_2/w_n133_n65#
+ VSUBS ypredec1_xa_3v1024x8m81_7/a_145_n4683# ypredec1_xa_3v1024x8m81_5/a_465_n4683#
+ ypredec1_xa_3v1024x8m81_7/a_0_56# ypredec1_xa_3v1024x8m81_7/a_465_n4683# ypredec1_xa_3v1024x8m81_6/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_3/a_145_n4683# ypredec1_xa_3v1024x8m81_7/a_305_n4683# ypredec1_xa_3v1024x8m81_7/a_305_n4683#
+ ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/pmos_5p04310591302060_3v1024x8m81_0/S
+ ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47821868_3v1024x8m81_3/w_n133_n66# ypredec1_xa_3v1024x8m81
.ends

.subckt ypredec1_bot_3v1024x8m81 pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ m1_n9_2295# m1_n9_2436# m1_n9_2154# m1_n9_2013# alatch_3v1024x8m81_0/a m3_10_2563#
+ m1_n9_1871# pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/S
+ m1_n9_1730# alatch_3v1024x8m81_0/enb VSUBS pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ alatch_3v1024x8m81_0/vdd
Xpmos_1p2$$46887980_3v1024x8m81_0 pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/S
+ pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/S pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D pmos_1p2$$46887980_3v1024x8m81
Xpmos_1p2$$46887980_3v1024x8m81_1 pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/S
+ pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/S pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ alatch_3v1024x8m81_0/ab pmos_1p2$$46887980_3v1024x8m81
Xalatch_3v1024x8m81_0 alatch_3v1024x8m81_0/en alatch_3v1024x8m81_0/ab alatch_3v1024x8m81_0/a
+ alatch_3v1024x8m81_0/vdd alatch_3v1024x8m81_0/enb m3_10_2563# VSUBS alatch_3v1024x8m81
Xnmos_1p2$$47514668_3v1024x8m81_0 VSUBS pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D VSUBS nmos_1p2$$47514668_3v1024x8m81
Xnmos_1p2$$47514668_3v1024x8m81_1 VSUBS pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ alatch_3v1024x8m81_0/ab VSUBS nmos_1p2$$47514668_3v1024x8m81
.ends

.subckt ypredec1_3v1024x8m81 ly[5] ly[4] ly[7] ly[3] ly[2] ly[1] ly[0] ry[0] ry[1]
+ ry[2] ry[3] ry[4] ry[5] ry[6] ry[7] ly[6] men A[0] A[1] A[2] clk ypredec1_bot_3v1024x8m81_0/alatch_3v1024x8m81_0/a
+ ypredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/a pmos_1p2$$47109164_3v1024x8m81_0/pmos_5p04310591302062_3v1024x8m81_0/S
+ ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/S
+ pmos_1p2$$47109164_3v1024x8m81_0/pmos_5p04310591302062_3v1024x8m81_0/w_n202_n86#
+ ypredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/vdd M1_NWELL13_3v1024x8m81_0/VSUBS
+ ypredec1_bot_3v1024x8m81_1/alatch_3v1024x8m81_0/a ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
Xypredec1_ys_3v1024x8m81_8 ry[6] ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ry[6] M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81
Xypredec1_ys_3v1024x8m81_9 ry[7] ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_3/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ry[7] M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81
Xnmos_1p2$$47342636_3v1024x8m81_0 M1_NWELL13_3v1024x8m81_0/VSUBS nmos_5p04310591302056_3v1024x8m81_1/D
+ ypredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/enb M1_NWELL13_3v1024x8m81_0/VSUBS
+ nmos_1p2$$47342636_3v1024x8m81
Xypredec1_ys_3v1024x8m81_10 ry[1] ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_1/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ry[1] M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81
Xypredec1_ys_3v1024x8m81_11 ry[2] ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_4/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ry[2] M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81
Xypredec1_ys_3v1024x8m81_12 ry[3] ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_0/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ry[3] M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81
Xypredec1_ys_3v1024x8m81_13 ry[4] ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_6/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ry[4] M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81
Xypredec1_ys_3v1024x8m81_14 ry[0] ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_5/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ry[0] M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81
Xypredec1_ys_3v1024x8m81_15 ly[7] ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_3/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ly[7] M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81
Xnmos_5p04310591302056_3v1024x8m81_0 M1_NWELL13_3v1024x8m81_0/VSUBS clk nmos_5p04310591302056_3v1024x8m81_1/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS nmos_5p04310591302056_3v1024x8m81
Xnmos_5p04310591302056_3v1024x8m81_1 nmos_5p04310591302056_3v1024x8m81_1/D men M1_NWELL13_3v1024x8m81_0/VSUBS
+ M1_NWELL13_3v1024x8m81_0/VSUBS nmos_5p04310591302056_3v1024x8m81
Xypredec1_xax8_3v1024x8m81_0 ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_6/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_5/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_3/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_4/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/S
+ ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_0/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_1/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_2/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_0/pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_1/pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_0/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/S
+ ypredec1_bot_3v1024x8m81_1/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/S
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_xax8_3v1024x8m81
Xpmos_1p2$$47109164_3v1024x8m81_0 pmos_1p2$$47109164_3v1024x8m81_0/pmos_5p04310591302062_3v1024x8m81_0/w_n202_n86#
+ ypredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/enb pmos_1p2$$47109164_3v1024x8m81_0/pmos_5p04310591302062_3v1024x8m81_0/S
+ nmos_5p04310591302056_3v1024x8m81_1/D pmos_1p2$$47109164_3v1024x8m81_0/pmos_5p04310591302062_3v1024x8m81_0/S
+ nmos_5p04310591302056_3v1024x8m81_1/D pmos_1p2$$47109164_3v1024x8m81
Xypredec1_ys_3v1024x8m81_0 ly[3] ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_0/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ly[3] M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81
Xypredec1_ys_3v1024x8m81_1 ly[4] ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_6/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ly[4] M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81
Xypredec1_ys_3v1024x8m81_2 ly[5] ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_2/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ly[5] M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81
Xypredec1_ys_3v1024x8m81_3 ly[6] ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_7/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ly[6] M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81
Xypredec1_ys_3v1024x8m81_4 ly[0] ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_5/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ly[0] M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81
Xypredec1_bot_3v1024x8m81_0 ypredec1_bot_3v1024x8m81_0/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_1/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_0/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_1/pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_0/alatch_3v1024x8m81_0/a nmos_5p04310591302056_3v1024x8m81_1/D
+ ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/S
+ ypredec1_bot_3v1024x8m81_0/pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/enb M1_NWELL13_3v1024x8m81_0/VSUBS
+ ypredec1_bot_3v1024x8m81_0/pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/vdd ypredec1_bot_3v1024x8m81
Xypredec1_bot_3v1024x8m81_1 ypredec1_bot_3v1024x8m81_1/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_1/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_0/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_1/pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_1/alatch_3v1024x8m81_0/a nmos_5p04310591302056_3v1024x8m81_1/D
+ ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/S
+ ypredec1_bot_3v1024x8m81_0/pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/enb M1_NWELL13_3v1024x8m81_0/VSUBS
+ ypredec1_bot_3v1024x8m81_1/pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/vdd ypredec1_bot_3v1024x8m81
Xypredec1_ys_3v1024x8m81_5 ly[1] ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_1/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ly[1] M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81
Xypredec1_bot_3v1024x8m81_2 ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_1/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_0/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_1/pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/a nmos_5p04310591302056_3v1024x8m81_1/D
+ ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_1/pmos_5p0431059130204_3v1024x8m81_0/S
+ ypredec1_bot_3v1024x8m81_0/pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/enb M1_NWELL13_3v1024x8m81_0/VSUBS
+ ypredec1_bot_3v1024x8m81_2/pmos_1p2$$46887980_3v1024x8m81_0/pmos_5p0431059130204_3v1024x8m81_0/D
+ ypredec1_bot_3v1024x8m81_2/alatch_3v1024x8m81_0/vdd ypredec1_bot_3v1024x8m81
Xypredec1_ys_3v1024x8m81_6 ly[2] ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_4/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ly[2] M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81
Xypredec1_ys_3v1024x8m81_7 ry[5] ypredec1_xax8_3v1024x8m81_0/ypredec1_xa_3v1024x8m81_2/pmos_1p2$$47820844_3v1024x8m81_2/pmos_5p04310591302061_3v1024x8m81_0/D
+ ry[5] M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81_9/pmos_5p04310591302055_3v1024x8m81_3/D
+ M1_NWELL13_3v1024x8m81_0/VSUBS ypredec1_ys_3v1024x8m81
X0 a_5490_186# clk nmos_5p04310591302056_3v1024x8m81_1/D pmos_1p2$$47109164_3v1024x8m81_0/pmos_5p04310591302062_3v1024x8m81_0/S pfet_03v3 ad=0.1917p pd=1.425u as=0.34345p ps=1.71u w=1.065u l=0.28u
X1 nmos_5p04310591302056_3v1024x8m81_1/D clk a_5176_186# pmos_1p2$$47109164_3v1024x8m81_0/pmos_5p04310591302062_3v1024x8m81_0/S pfet_03v3 ad=0.34345p pd=1.71u as=0.19435p ps=1.43u w=1.065u l=0.28u
X2 a_5176_186# men pmos_1p2$$47109164_3v1024x8m81_0/pmos_5p04310591302062_3v1024x8m81_0/S pmos_1p2$$47109164_3v1024x8m81_0/pmos_5p04310591302062_3v1024x8m81_0/S pfet_03v3 ad=0.19435p pd=1.43u as=0.59108p ps=3.24u w=1.065u l=0.28u
X3 pmos_1p2$$47109164_3v1024x8m81_0/pmos_5p04310591302062_3v1024x8m81_0/S men a_5490_186# pmos_1p2$$47109164_3v1024x8m81_0/pmos_5p04310591302062_3v1024x8m81_0/S pfet_03v3 ad=0.59108p pd=3.24u as=0.1917p ps=1.425u w=1.065u l=0.28u
.ends

.subckt control_3v1024x8_3v1024x8m81 RYS[7] RYS[6] RYS[5] RYS[4] RYS[3] RYS[2] RYS[1]
+ RYS[0] LYS[0] LYS[1] LYS[2] LYS[3] LYS[6] LYS[5] LYS[4] LYS[7] tblhl IGWEN xb[3]
+ xb[2] xb[0] xa[7] xa[6] xa[5] xa[4] xa[2] A[0] xb[1] xc[3] xc[2] xa[1] A[9] A[7]
+ CLK A[2] A[1] A[6] A[3] A[4] A[5] A[8] GWEN VDD_uq0 VDD_uq5 VDD_uq6 VSS_uq2 VDD_uq4
+ xa[0] xa[3] men CEN gen_3v1024x8_3v1024x8m81_0/VDD_uq2 xc[1] VDD xc[0] GWE VDD_uq1
+ VDD_uq2 VSS
Xprexdec_top_3v1024x8m81_0 A[9] A[7] xb[3] xc[2] xb[1] xb[2] xb[0] xa[1] xa[2] xa[4]
+ xa[5] xa[6] xa[7] A[3] A[6] A[8] A[4] CLK VDD VDD xa[0] A[5] xa[3] xc[1] xc[0] VDD_uq1
+ men xc[3] VDD_uq1 CLK VSS VDD prexdec_top_3v1024x8m81
Xgen_3v1024x8_3v1024x8m81_0 VSS tblhl CEN CLK gen_3v1024x8_3v1024x8m81_0/WEN GWE GWEN
+ VDD_uq2 VDD_uq4 men gen_3v1024x8_3v1024x8m81_0/pmos_5p04310591302088_3v1024x8m81_0/D
+ IGWEN gen_3v1024x8_3v1024x8m81_0/VDD_uq2 gen_3v1024x8_3v1024x8m81
Xypredec1_3v1024x8m81_0 LYS[5] LYS[4] LYS[7] LYS[3] LYS[2] LYS[1] LYS[0] RYS[0] RYS[1]
+ RYS[2] RYS[3] RYS[4] RYS[5] RYS[6] RYS[7] LYS[6] men A[0] A[1] A[2] CLK A[0] A[1]
+ VDD_uq4 VDD_uq6 VDD_uq4 VDD_uq5 VSS A[2] VDD_uq2 ypredec1_3v1024x8m81
.ends

.subckt pmos_5p043105913020104_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.4004p pd=2.06u as=0.6776p ps=3.96u w=1.54u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.6776p pd=3.96u as=0.4004p ps=2.06u w=1.54u l=0.28u
.ends

.subckt pmos_1p2_02_R270_3v1024x8m81 a_118_n33# a_n41_n33# pmos_5p043105913020104_3v1024x8m81_0/S_uq0
+ w_n138_n63# pmos_5p043105913020104_3v1024x8m81_0/S pmos_5p043105913020104_3v1024x8m81_0/D
Xpmos_5p043105913020104_3v1024x8m81_0 pmos_5p043105913020104_3v1024x8m81_0/D a_n41_n33#
+ a_118_n33# w_n138_n63# pmos_5p043105913020104_3v1024x8m81_0/S_uq0 pmos_5p043105913020104_3v1024x8m81_0/S
+ pmos_5p043105913020104_3v1024x8m81
.ends

.subckt pmos_5p043105913020108_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.6669p pd=3.085u as=1.1286p ps=6.01u w=2.565u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=1.1286p pd=6.01u as=0.6669p ps=3.085u w=2.565u l=0.28u
.ends

.subckt pmos_1p2_01_R270_3v1024x8m81 pmos_5p043105913020108_3v1024x8m81_0/D w_n246_n93#
+ pmos_5p043105913020108_3v1024x8m81_0/S_uq0 pmos_5p043105913020108_3v1024x8m81_0/S
+ a_118_n33# a_n41_n33#
Xpmos_5p043105913020108_3v1024x8m81_0 pmos_5p043105913020108_3v1024x8m81_0/D a_n41_n33#
+ a_118_n33# w_n246_n93# pmos_5p043105913020108_3v1024x8m81_0/S_uq0 pmos_5p043105913020108_3v1024x8m81_0/S
+ pmos_5p043105913020108_3v1024x8m81
.ends

.subckt nmos_5p043105913020107_3v1024x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.6058p pd=2.85u as=1.0252p ps=5.54u w=2.33u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=1.0252p pd=5.54u as=0.6058p ps=2.85u w=2.33u l=0.28u
.ends

.subckt pmos_5p043105913020110_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.3256p pd=2.36u as=0.3256p ps=2.36u w=0.74u l=0.28u
.ends

.subckt nmos_5p043105913020109_3v1024x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.4004p pd=2.06u as=0.6776p ps=3.96u w=1.54u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.6776p pd=3.96u as=0.4004p ps=2.06u w=1.54u l=0.28u
.ends

.subckt pmos_5p043105913020103_3v1024x8m81 D_uq0 D a_265_n44# S_uq0 S a_n56_n44# a_104_n44#
+ w_n230_n86#
X0 D_uq0 a_265_n44# S_uq0 w_n230_n86# pfet_03v3 ad=2.0526p pd=10.21u as=1.22455p ps=5.19u w=4.665u l=0.28u
X1 D a_n56_n44# S w_n230_n86# pfet_03v3 ad=1.2129p pd=5.185u as=2.0526p ps=10.21u w=4.665u l=0.28u
X2 S_uq0 a_104_n44# D w_n230_n86# pfet_03v3 ad=1.22455p pd=5.19u as=1.2129p ps=5.185u w=4.665u l=0.28u
.ends

.subckt nmos_5p043105913020106_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1601p pd=1.64u as=0.1601p ps=1.64u w=0.305u l=0.28u
.ends

.subckt nmos_1p2_02_R270_3v1024x8m81 nmos_5p04310591302044_3v1024x8m81_0/D a_n14_n33#
+ VSUBS nmos_5p04310591302044_3v1024x8m81_0/S
Xnmos_5p04310591302044_3v1024x8m81_0 nmos_5p04310591302044_3v1024x8m81_0/D a_n14_n33#
+ nmos_5p04310591302044_3v1024x8m81_0/S VSUBS nmos_5p04310591302044_3v1024x8m81
.ends

.subckt pmos_5p043105913020105_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.28u
.ends

.subckt pmos_1p2_03_R270_3v1024x8m81 pmos_5p043105913020103_3v1024x8m81_0/D_uq0 pmos_5p043105913020103_3v1024x8m81_0/D
+ a_n69_n138# w_n138_n63# pmos_5p043105913020103_3v1024x8m81_0/S_uq0 a_90_n138# pmos_5p043105913020103_3v1024x8m81_0/S
+ a_251_n138#
Xpmos_5p043105913020103_3v1024x8m81_0 pmos_5p043105913020103_3v1024x8m81_0/D_uq0 pmos_5p043105913020103_3v1024x8m81_0/D
+ a_251_n138# pmos_5p043105913020103_3v1024x8m81_0/S_uq0 pmos_5p043105913020103_3v1024x8m81_0/S
+ a_n69_n138# a_90_n138# w_n138_n63# pmos_5p043105913020103_3v1024x8m81
.ends

.subckt xdec_3v1024x8m81 RWL LWL men xc xb xa m2_11898_n156# m2_9070_n156# m2_7748_n156#
+ m2_8806_n156# m2_10577_n156# m2_10840_n156# m2_7219_n156# m2_7483_n156# m2_11634_n156#
+ m2_8277_n156# m2_12427_n156# m2_8541_n156# m2_11105_n156# m2_11370_n156# m2_8012_n156#
+ m2_12163_n156# vdd vss
Xpmos_1p2_02_R270_3v1024x8m81_0 pmos_5p043105913020105_3v1024x8m81_3/S pmos_5p043105913020105_3v1024x8m81_3/S
+ nmos_5p043105913020109_3v1024x8m81_0/S vdd nmos_5p043105913020109_3v1024x8m81_0/S
+ men pmos_1p2_02_R270_3v1024x8m81
Xpmos_1p2_01_R270_3v1024x8m81_0 pmos_1p2_01_R270_3v1024x8m81_0/pmos_5p043105913020108_3v1024x8m81_0/D
+ vdd vdd vdd nmos_5p043105913020109_3v1024x8m81_0/S nmos_5p043105913020109_3v1024x8m81_0/S
+ pmos_1p2_01_R270_3v1024x8m81
Xpmos_1p2_01_R270_3v1024x8m81_1 pmos_1p2_01_R270_3v1024x8m81_1/pmos_5p043105913020108_3v1024x8m81_0/D
+ vdd vdd vdd nmos_5p043105913020109_3v1024x8m81_0/S nmos_5p043105913020109_3v1024x8m81_0/S
+ pmos_1p2_01_R270_3v1024x8m81
Xnmos_5p043105913020107_3v1024x8m81_0 LWL pmos_1p2_01_R270_3v1024x8m81_1/pmos_5p043105913020108_3v1024x8m81_0/D
+ pmos_1p2_01_R270_3v1024x8m81_1/pmos_5p043105913020108_3v1024x8m81_0/D vss vss vss
+ nmos_5p043105913020107_3v1024x8m81
Xnmos_5p043105913020107_3v1024x8m81_1 RWL pmos_1p2_01_R270_3v1024x8m81_0/pmos_5p043105913020108_3v1024x8m81_0/D
+ pmos_1p2_01_R270_3v1024x8m81_0/pmos_5p043105913020108_3v1024x8m81_0/D vss vss vss
+ nmos_5p043105913020107_3v1024x8m81
Xpmos_5p043105913020110_3v1024x8m81_0 vdd pmos_5p043105913020105_3v1024x8m81_3/S vdd
+ pmos_5p043105913020110_3v1024x8m81_0/S pmos_5p043105913020110_3v1024x8m81
Xnmos_5p043105913020109_3v1024x8m81_0 men pmos_5p043105913020110_3v1024x8m81_0/S pmos_5p043105913020110_3v1024x8m81_0/S
+ nmos_5p043105913020109_3v1024x8m81_0/S nmos_5p043105913020109_3v1024x8m81_0/S vss
+ nmos_5p043105913020109_3v1024x8m81
Xpmos_5p043105913020103_3v1024x8m81_0 vdd vdd pmos_1p2_01_R270_3v1024x8m81_0/pmos_5p043105913020108_3v1024x8m81_0/D
+ RWL RWL pmos_1p2_01_R270_3v1024x8m81_0/pmos_5p043105913020108_3v1024x8m81_0/D pmos_1p2_01_R270_3v1024x8m81_0/pmos_5p043105913020108_3v1024x8m81_0/D
+ vdd pmos_5p043105913020103_3v1024x8m81
Xnmos_5p043105913020106_3v1024x8m81_0 vss pmos_5p043105913020105_3v1024x8m81_3/S pmos_5p043105913020110_3v1024x8m81_0/S
+ vss nmos_5p043105913020106_3v1024x8m81
Xnmos_1p2_02_R270_3v1024x8m81_0 vss pmos_5p043105913020105_3v1024x8m81_3/S vss nmos_5p043105913020109_3v1024x8m81_0/S
+ nmos_1p2_02_R270_3v1024x8m81
Xpmos_5p043105913020105_3v1024x8m81_1 pmos_5p043105913020105_3v1024x8m81_3/S xb vdd
+ vdd pmos_5p043105913020105_3v1024x8m81
Xpmos_5p043105913020105_3v1024x8m81_2 vdd xa vdd pmos_5p043105913020105_3v1024x8m81_3/S
+ pmos_5p043105913020105_3v1024x8m81
Xpmos_5p043105913020105_3v1024x8m81_3 vdd xc vdd pmos_5p043105913020105_3v1024x8m81_3/S
+ pmos_5p043105913020105_3v1024x8m81
Xpmos_1p2_03_R270_3v1024x8m81_0 vdd vdd pmos_1p2_01_R270_3v1024x8m81_1/pmos_5p043105913020108_3v1024x8m81_0/D
+ vdd LWL pmos_1p2_01_R270_3v1024x8m81_1/pmos_5p043105913020108_3v1024x8m81_0/D LWL
+ pmos_1p2_01_R270_3v1024x8m81_1/pmos_5p043105913020108_3v1024x8m81_0/D pmos_1p2_03_R270_3v1024x8m81
X0 vss xc a_9450_422# vss nfet_03v3 ad=0.88935p pd=4.15u as=0.29032p ps=1.865u w=1.47u l=0.28u
X1 vss nmos_5p043105913020109_3v1024x8m81_0/S pmos_1p2_01_R270_3v1024x8m81_1/pmos_5p043105913020108_3v1024x8m81_0/D vss nfet_03v3 ad=0.2796p pd=4.9u as=1.0252p ps=5.54u w=2.33u l=0.28u
X2 a_9450_280# xa pmos_5p043105913020105_3v1024x8m81_3/S vss nfet_03v3 ad=0.31605p pd=1.9u as=0.74235p ps=3.95u w=1.47u l=0.28u
X3 a_9450_422# xb a_9450_280# vss nfet_03v3 ad=0.29032p pd=1.865u as=0.31605p ps=1.9u w=1.47u l=0.28u
X4 vss nmos_5p043105913020109_3v1024x8m81_0/S pmos_1p2_01_R270_3v1024x8m81_0/pmos_5p043105913020108_3v1024x8m81_0/D vss nfet_03v3 ad=1.15335p pd=5.65u as=1.0718p ps=5.58u w=2.33u l=0.28u
.ends

.subckt xdec8_3v1024x8m81 LWL[4] LWL[2] RWL[5] RWL[2] RWL[6] LWL[1] LWL[7] LWL[6]
+ LWL[0] LWL[3] RWL[3] xc xb xa[4] xa[7] xb_uq3 xc_uq0 xc_uq2 xc_uq3 xc_uq6 xb_uq6
+ xa[1] xdec_3v1024x8m81_7/m2_12163_n156# RWL[0] xb_uq2 xc_uq5 xdec_3v1024x8m81_7/m2_8806_n156#
+ xb_uq0 xa[3] xb_uq5 xa[0] xa[6] xdec_3v1024x8m81_7/m2_10577_n156# RWL[1] xdec_3v1024x8m81_7/m2_10840_n156#
+ xdec_3v1024x8m81_7/m2_8277_n156# xdec_3v1024x8m81_7/m2_8012_n156# RWL[7] LWL[5]
+ xc_uq4 xc_uq1 xb_uq4 xdec_3v1024x8m81_7/m2_11634_n156# xdec_3v1024x8m81_7/m2_8541_n156#
+ RWL[4] xb_uq1 xdec_3v1024x8m81_7/m2_11105_n156# xa[5] xdec_3v1024x8m81_7/m2_7219_n156#
+ xa[2] xdec_3v1024x8m81_7/m2_12427_n156# xdec_3v1024x8m81_7/m2_7483_n156# men xdec_3v1024x8m81_7/m2_9070_n156#
+ xdec_3v1024x8m81_7/m2_7748_n156# xdec_3v1024x8m81_7/m2_11898_n156# xdec_3v1024x8m81_7/m2_11370_n156#
+ vdd vss
Xxdec_3v1024x8m81_0 RWL[6] LWL[6] men xc_uq5 xb_uq5 xa[6] xdec_3v1024x8m81_7/m2_11898_n156#
+ xdec_3v1024x8m81_7/m2_9070_n156# xdec_3v1024x8m81_7/m2_7748_n156# xdec_3v1024x8m81_7/m2_8806_n156#
+ xdec_3v1024x8m81_7/m2_10577_n156# xdec_3v1024x8m81_7/m2_10840_n156# xdec_3v1024x8m81_7/m2_7219_n156#
+ xdec_3v1024x8m81_7/m2_7483_n156# xdec_3v1024x8m81_7/m2_11634_n156# xdec_3v1024x8m81_7/m2_8277_n156#
+ xdec_3v1024x8m81_7/m2_12427_n156# xdec_3v1024x8m81_7/m2_8541_n156# xdec_3v1024x8m81_7/m2_11105_n156#
+ xdec_3v1024x8m81_7/m2_11370_n156# xdec_3v1024x8m81_7/m2_8012_n156# xdec_3v1024x8m81_7/m2_12163_n156#
+ vdd vss xdec_3v1024x8m81
Xxdec_3v1024x8m81_1 RWL[4] LWL[4] men xc_uq3 xb_uq3 xa[4] xdec_3v1024x8m81_7/m2_11898_n156#
+ xdec_3v1024x8m81_7/m2_9070_n156# xdec_3v1024x8m81_7/m2_7748_n156# xdec_3v1024x8m81_7/m2_8806_n156#
+ xdec_3v1024x8m81_7/m2_10577_n156# xdec_3v1024x8m81_7/m2_10840_n156# xdec_3v1024x8m81_7/m2_7219_n156#
+ xdec_3v1024x8m81_7/m2_7483_n156# xdec_3v1024x8m81_7/m2_11634_n156# xdec_3v1024x8m81_7/m2_8277_n156#
+ xdec_3v1024x8m81_7/m2_12427_n156# xdec_3v1024x8m81_7/m2_8541_n156# xdec_3v1024x8m81_7/m2_11105_n156#
+ xdec_3v1024x8m81_7/m2_11370_n156# xdec_3v1024x8m81_7/m2_8012_n156# xdec_3v1024x8m81_7/m2_12163_n156#
+ vdd vss xdec_3v1024x8m81
Xxdec_3v1024x8m81_2 RWL[2] LWL[2] men xc_uq1 xb_uq1 xa[2] xdec_3v1024x8m81_7/m2_11898_n156#
+ xdec_3v1024x8m81_7/m2_9070_n156# xdec_3v1024x8m81_7/m2_7748_n156# xdec_3v1024x8m81_7/m2_8806_n156#
+ xdec_3v1024x8m81_7/m2_10577_n156# xdec_3v1024x8m81_7/m2_10840_n156# xdec_3v1024x8m81_7/m2_7219_n156#
+ xdec_3v1024x8m81_7/m2_7483_n156# xdec_3v1024x8m81_7/m2_11634_n156# xdec_3v1024x8m81_7/m2_8277_n156#
+ xdec_3v1024x8m81_7/m2_12427_n156# xdec_3v1024x8m81_7/m2_8541_n156# xdec_3v1024x8m81_7/m2_11105_n156#
+ xdec_3v1024x8m81_7/m2_11370_n156# xdec_3v1024x8m81_7/m2_8012_n156# xdec_3v1024x8m81_7/m2_12163_n156#
+ vdd vss xdec_3v1024x8m81
Xxdec_3v1024x8m81_3 RWL[0] LWL[0] men xc_uq0 xb_uq0 xa[0] xdec_3v1024x8m81_7/m2_11898_n156#
+ xdec_3v1024x8m81_7/m2_9070_n156# xdec_3v1024x8m81_7/m2_7748_n156# xdec_3v1024x8m81_7/m2_8806_n156#
+ xdec_3v1024x8m81_7/m2_10577_n156# xdec_3v1024x8m81_7/m2_10840_n156# xdec_3v1024x8m81_7/m2_7219_n156#
+ xdec_3v1024x8m81_7/m2_7483_n156# xdec_3v1024x8m81_7/m2_11634_n156# xdec_3v1024x8m81_7/m2_8277_n156#
+ xdec_3v1024x8m81_7/m2_12427_n156# xdec_3v1024x8m81_7/m2_8541_n156# xdec_3v1024x8m81_7/m2_11105_n156#
+ xdec_3v1024x8m81_7/m2_11370_n156# xdec_3v1024x8m81_7/m2_8012_n156# xdec_3v1024x8m81_7/m2_12163_n156#
+ vdd vss xdec_3v1024x8m81
Xxdec_3v1024x8m81_4 RWL[7] LWL[7] men xc_uq6 xb_uq6 xa[7] xdec_3v1024x8m81_7/m2_11898_n156#
+ xdec_3v1024x8m81_7/m2_9070_n156# xdec_3v1024x8m81_7/m2_7748_n156# xdec_3v1024x8m81_7/m2_8806_n156#
+ xdec_3v1024x8m81_7/m2_10577_n156# xdec_3v1024x8m81_7/m2_10840_n156# xdec_3v1024x8m81_7/m2_7219_n156#
+ xdec_3v1024x8m81_7/m2_7483_n156# xdec_3v1024x8m81_7/m2_11634_n156# xdec_3v1024x8m81_7/m2_8277_n156#
+ xdec_3v1024x8m81_7/m2_12427_n156# xdec_3v1024x8m81_7/m2_8541_n156# xdec_3v1024x8m81_7/m2_11105_n156#
+ xdec_3v1024x8m81_7/m2_11370_n156# xdec_3v1024x8m81_7/m2_8012_n156# xdec_3v1024x8m81_7/m2_12163_n156#
+ vdd vss xdec_3v1024x8m81
Xxdec_3v1024x8m81_5 RWL[5] LWL[5] men xc_uq4 xb_uq4 xa[5] xdec_3v1024x8m81_7/m2_11898_n156#
+ xdec_3v1024x8m81_7/m2_9070_n156# xdec_3v1024x8m81_7/m2_7748_n156# xdec_3v1024x8m81_7/m2_8806_n156#
+ xdec_3v1024x8m81_7/m2_10577_n156# xdec_3v1024x8m81_7/m2_10840_n156# xdec_3v1024x8m81_7/m2_7219_n156#
+ xdec_3v1024x8m81_7/m2_7483_n156# xdec_3v1024x8m81_7/m2_11634_n156# xdec_3v1024x8m81_7/m2_8277_n156#
+ xdec_3v1024x8m81_7/m2_12427_n156# xdec_3v1024x8m81_7/m2_8541_n156# xdec_3v1024x8m81_7/m2_11105_n156#
+ xdec_3v1024x8m81_7/m2_11370_n156# xdec_3v1024x8m81_7/m2_8012_n156# xdec_3v1024x8m81_7/m2_12163_n156#
+ vdd vss xdec_3v1024x8m81
Xxdec_3v1024x8m81_6 RWL[3] LWL[3] men xc_uq2 xb_uq2 xa[3] xdec_3v1024x8m81_7/m2_11898_n156#
+ xdec_3v1024x8m81_7/m2_9070_n156# xdec_3v1024x8m81_7/m2_7748_n156# xdec_3v1024x8m81_7/m2_8806_n156#
+ xdec_3v1024x8m81_7/m2_10577_n156# xdec_3v1024x8m81_7/m2_10840_n156# xdec_3v1024x8m81_7/m2_7219_n156#
+ xdec_3v1024x8m81_7/m2_7483_n156# xdec_3v1024x8m81_7/m2_11634_n156# xdec_3v1024x8m81_7/m2_8277_n156#
+ xdec_3v1024x8m81_7/m2_12427_n156# xdec_3v1024x8m81_7/m2_8541_n156# xdec_3v1024x8m81_7/m2_11105_n156#
+ xdec_3v1024x8m81_7/m2_11370_n156# xdec_3v1024x8m81_7/m2_8012_n156# xdec_3v1024x8m81_7/m2_12163_n156#
+ vdd vss xdec_3v1024x8m81
Xxdec_3v1024x8m81_7 RWL[1] LWL[1] men xc xb xa[1] xdec_3v1024x8m81_7/m2_11898_n156#
+ xdec_3v1024x8m81_7/m2_9070_n156# xdec_3v1024x8m81_7/m2_7748_n156# xdec_3v1024x8m81_7/m2_8806_n156#
+ xdec_3v1024x8m81_7/m2_10577_n156# xdec_3v1024x8m81_7/m2_10840_n156# xdec_3v1024x8m81_7/m2_7219_n156#
+ xdec_3v1024x8m81_7/m2_7483_n156# xdec_3v1024x8m81_7/m2_11634_n156# xdec_3v1024x8m81_7/m2_8277_n156#
+ xdec_3v1024x8m81_7/m2_12427_n156# xdec_3v1024x8m81_7/m2_8541_n156# xdec_3v1024x8m81_7/m2_11105_n156#
+ xdec_3v1024x8m81_7/m2_11370_n156# xdec_3v1024x8m81_7/m2_8012_n156# xdec_3v1024x8m81_7/m2_12163_n156#
+ vdd vss xdec_3v1024x8m81
.ends

.subckt xdec64_468_3v1024x8m81 LWL[6] LWL[7] RWL[18] RWL[17] RWL[15] RWL[14] RWL[13]
+ LWL[9] LWL[8] LWL[0] LWL[1] LWL[2] LWL[3] LWL[4] LWL[5] RWL[11] RWL[10] RWL[9] RWL[8]
+ RWL[7] RWL[5] RWL[1] RWL[0] LWL[18] LWL[17] LWL[16] LWL[15] LWL[14] LWL[13] LWL[12]
+ LWL[11] LWL[10] RWL[4] LWL[28] LWL[27] LWL[26] LWL[25] LWL[24] LWL[23] LWL[22] LWL[21]
+ LWL[20] LWL[19] RWL[22] RWL[26] RWL[27] RWL[30] RWL[31] LWL[31] LWL[30] LWL[29]
+ xa[0] xa[3] xa[4] xa[5] xa[6] xa[7] xb[3] xb[2] xb[1] xb[0] xc xa[1] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_8012_n156#
+ RWL[23] RWL[20] RWL[24] RWL[21] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7483_n156#
+ xa[2] RWL[2] RWL[25] RWL[28] RWL[12] RWL[3] men RWL[19] xdec8_3v1024x8m81_3/xc RWL[16]
+ RWL[6] RWL[29] vdd vss
Xxdec8_3v1024x8m81_0 LWL[28] LWL[26] RWL[29] RWL[26] RWL[30] LWL[25] LWL[31] LWL[30]
+ LWL[24] LWL[27] RWL[27] xdec8_3v1024x8m81_3/xc xb[3] xa[4] xa[7] xb[3] xdec8_3v1024x8m81_3/xc
+ xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xb[3] xa[1]
+ xa[1] RWL[24] xb[3] xdec8_3v1024x8m81_3/xc xb[1] xb[3] xa[3] xb[3] xa[0] xa[6] xa[7]
+ RWL[25] xa[6] xb[3] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_8012_n156# RWL[31]
+ LWL[29] xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xb[3] xa[3] xb[2] RWL[28]
+ xb[3] xa[5] xa[5] xdec8_3v1024x8m81_3/xc xa[2] xa[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7483_n156#
+ men xb[0] xc xa[2] xa[4] vdd vss xdec8_3v1024x8m81
Xxdec8_3v1024x8m81_1 LWL[4] LWL[2] RWL[5] RWL[2] RWL[6] LWL[1] LWL[7] LWL[6] LWL[0]
+ LWL[3] RWL[3] xdec8_3v1024x8m81_3/xc xb[0] xa[4] xa[7] xb[0] xdec8_3v1024x8m81_3/xc
+ xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xb[0] xa[1]
+ xa[1] RWL[0] xb[0] xdec8_3v1024x8m81_3/xc xb[1] xb[0] xa[3] xb[0] xa[0] xa[6] xa[7]
+ RWL[1] xa[6] xb[3] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_8012_n156# RWL[7] LWL[5]
+ xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xb[0] xa[3] xb[2] RWL[4] xb[0] xa[5]
+ xa[5] xdec8_3v1024x8m81_3/xc xa[2] xa[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7483_n156#
+ men xb[0] xc xa[2] xa[4] vdd vss xdec8_3v1024x8m81
Xxdec8_3v1024x8m81_2 LWL[12] LWL[10] RWL[13] RWL[10] RWL[14] LWL[9] LWL[15] LWL[14]
+ LWL[8] LWL[11] RWL[11] xdec8_3v1024x8m81_3/xc xb[1] xa[4] xa[7] xb[1] xdec8_3v1024x8m81_3/xc
+ xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xb[1] xa[1]
+ xa[1] RWL[8] xb[1] xdec8_3v1024x8m81_3/xc xb[1] xb[1] xa[3] xb[1] xa[0] xa[6] xa[7]
+ RWL[9] xa[6] xb[3] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_8012_n156# RWL[15]
+ LWL[13] xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xb[1] xa[3] xb[2] RWL[12]
+ xb[1] xa[5] xa[5] xdec8_3v1024x8m81_3/xc xa[2] xa[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7483_n156#
+ men xb[0] xc xa[2] xa[4] vdd vss xdec8_3v1024x8m81
Xxdec8_3v1024x8m81_3 LWL[20] LWL[18] RWL[21] RWL[18] RWL[22] LWL[17] LWL[23] LWL[22]
+ LWL[16] LWL[19] RWL[19] xdec8_3v1024x8m81_3/xc xb[2] xa[4] xa[7] xb[2] xdec8_3v1024x8m81_3/xc
+ xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xb[2] xa[1]
+ xa[1] RWL[16] xb[2] xdec8_3v1024x8m81_3/xc xb[1] xb[2] xa[3] xb[2] xa[0] xa[6] xa[7]
+ RWL[17] xa[6] xb[3] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_8012_n156# RWL[23]
+ LWL[21] xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xb[2] xa[3] xb[2] RWL[20]
+ xb[2] xa[5] xa[5] xdec8_3v1024x8m81_3/xc xa[2] xa[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7483_n156#
+ men xb[0] xc xa[2] xa[4] vdd vss xdec8_3v1024x8m81
.ends

.subckt nmos_5p043105913020111_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.5412p pd=3.34u as=0.5412p ps=3.34u w=1.23u l=0.28u
.ends

.subckt pmos_5p043105913020101_3v1024x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=1.353p pd=7.03u as=1.353p ps=7.03u w=3.075u l=0.28u
.ends

.subckt pmos_1p2_01_R90_3v1024x8m81 pmos_5p043105913020101_3v1024x8m81_0/S w_n137_n63#
+ a_n14_n33# pmos_5p043105913020101_3v1024x8m81_0/D
Xpmos_5p043105913020101_3v1024x8m81_0 pmos_5p043105913020101_3v1024x8m81_0/D a_n14_n33#
+ w_n137_n63# pmos_5p043105913020101_3v1024x8m81_0/S pmos_5p043105913020101_3v1024x8m81
.ends

.subckt nmos_5p04310591302099_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=2.0746p pd=10.31u as=2.0746p ps=10.31u w=4.715u l=0.28u
.ends

.subckt nmos_1p2_02_R90_3v1024x8m81 nmos_5p04310591302099_3v1024x8m81_0/S nmos_5p04310591302099_3v1024x8m81_0/D
+ a_n14_n33# VSUBS
Xnmos_5p04310591302099_3v1024x8m81_0 nmos_5p04310591302099_3v1024x8m81_0/D a_n14_n33#
+ nmos_5p04310591302099_3v1024x8m81_0/S VSUBS nmos_5p04310591302099_3v1024x8m81
.ends

.subckt pmoscap_R270_3v1024x8m81 m3_770_16# a_n126_928# a_n140_236# m3_152_0# w_n226_n219#
X0 a_n140_236# a_n126_928# a_n140_236# w_n226_n219# pfet_03v3 ad=1.20555p pd=6.07u as=0 ps=0 w=2.565u l=2.505u
X1 a_n140_236# a_n126_928# a_n140_236# w_n226_n219# pfet_03v3 ad=0.6733p pd=3.09u as=0 ps=0 w=2.565u l=2.505u
.ends

.subckt xdec32_3v1024x8m81 LWL[6] LWL[7] RWL[18] RWL[17] RWL[15] RWL[14] RWL[13] LWL[9]
+ LWL[8] LWL[0] LWL[1] LWL[2] LWL[3] LWL[4] LWL[5] RWL[11] RWL[10] RWL[9] RWL[8] RWL[7]
+ RWL[5] RWL[1] LWL[18] LWL[17] LWL[16] LWL[15] LWL[14] LWL[13] LWL[12] LWL[11] LWL[10]
+ RWL[4] LWL[28] LWL[27] LWL[26] LWL[25] LWL[24] LWL[23] LWL[22] LWL[21] LWL[20] LWL[19]
+ RWL[22] RWL[23] RWL[26] RWL[27] RWL[30] RWL[31] LWL[31] LWL[30] LWL[29] xb[3] xb[2]
+ xb[1] xb[0] RWL[20] RWL[24] xa[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7219_n156#
+ RWL[21] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7483_n156# RWL[2] RWL[25] xc xa[5]
+ xa[4] RWL[28] RWL[12] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7748_n156# RWL[3]
+ men xa[1] xa[7] RWL[19] RWL[0] xa[6] RWL[16] xa[2] RWL[6] vdd RWL[29] xa[3] vss
Xxdec8_3v1024x8m81_0 LWL[28] LWL[26] RWL[29] RWL[26] RWL[30] LWL[25] LWL[31] LWL[30]
+ LWL[24] LWL[27] RWL[27] xc xb[3] xa[4] xa[7] xb[3] xc xc xc xc xb[3] xa[1] xa[1]
+ RWL[24] xb[3] xc xb[1] xb[3] xa[3] xb[3] xa[0] xa[6] xa[7] RWL[25] xa[6] xb[3] xc
+ RWL[31] LWL[29] xc xc xb[3] xa[3] xb[2] RWL[28] xb[3] xa[5] xa[5] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7219_n156#
+ xa[2] xa[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7483_n156# men xb[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7748_n156#
+ xa[2] xa[4] vdd vss xdec8_3v1024x8m81
Xxdec8_3v1024x8m81_1 LWL[4] LWL[2] RWL[5] RWL[2] RWL[6] LWL[1] LWL[7] LWL[6] LWL[0]
+ LWL[3] RWL[3] xc xb[0] xa[4] xa[7] xb[0] xc xc xc xc xb[0] xa[1] xa[1] RWL[0] xb[0]
+ xc xb[1] xb[0] xa[3] xb[0] xa[0] xa[6] xa[7] RWL[1] xa[6] xb[3] xc RWL[7] LWL[5]
+ xc xc xb[0] xa[3] xb[2] RWL[4] xb[0] xa[5] xa[5] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7219_n156#
+ xa[2] xa[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7483_n156# men xb[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7748_n156#
+ xa[2] xa[4] vdd vss xdec8_3v1024x8m81
Xxdec8_3v1024x8m81_2 LWL[12] LWL[10] RWL[13] RWL[10] RWL[14] LWL[9] LWL[15] LWL[14]
+ LWL[8] LWL[11] RWL[11] xc xb[1] xa[4] xa[7] xb[1] xc xc xc xc xb[1] xa[1] xa[1]
+ RWL[8] xb[1] xc xb[1] xb[1] xa[3] xb[1] xa[0] xa[6] xa[7] RWL[9] xa[6] xb[3] xc
+ RWL[15] LWL[13] xc xc xb[1] xa[3] xb[2] RWL[12] xb[1] xa[5] xa[5] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7219_n156#
+ xa[2] xa[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7483_n156# men xb[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7748_n156#
+ xa[2] xa[4] vdd vss xdec8_3v1024x8m81
Xxdec8_3v1024x8m81_3 LWL[20] LWL[18] RWL[21] RWL[18] RWL[22] LWL[17] LWL[23] LWL[22]
+ LWL[16] LWL[19] RWL[19] xc xb[2] xa[4] xa[7] xb[2] xc xc xc xc xb[2] xa[1] xa[1]
+ RWL[16] xb[2] xc xb[1] xb[2] xa[3] xb[2] xa[0] xa[6] xa[7] RWL[17] xa[6] xb[3] xc
+ RWL[23] LWL[21] xc xc xb[2] xa[3] xb[2] RWL[20] xb[2] xa[5] xa[5] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7219_n156#
+ xa[2] xa[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7483_n156# men xb[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7748_n156#
+ xa[2] xa[4] vdd vss xdec8_3v1024x8m81
.ends

.subckt pmoscap_L1_W2_R270_3v1024x8m81 m3_307_0# m3_600_0# M2_M1$04_R270_3v1024x8m81_0/VSUBS
+ a_597_236# a_8_236# m1_38_36#
X0 a_597_236# M2_M1$04_R270_3v1024x8m81_0/VSUBS a_8_236# m1_38_36# pfet_03v3 ad=1.1286p pd=6.01u as=1.1286p ps=6.01u w=2.565u l=2.505u
.ends

.subckt pmos_5p043105913020100_3v1024x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=1.5314p pd=6.41u as=2.5916p ps=12.66u w=5.89u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=2.5916p pd=12.66u as=1.5314p ps=6.41u w=5.89u l=0.28u
.ends

.subckt pmos_1p2_02_R90_3v1024x8m81 pmos_5p043105913020100_3v1024x8m81_0/S_uq0 pmos_5p043105913020100_3v1024x8m81_0/S
+ w_n138_n63# a_118_n33# pmos_5p043105913020100_3v1024x8m81_0/D a_n41_n33#
Xpmos_5p043105913020100_3v1024x8m81_0 pmos_5p043105913020100_3v1024x8m81_0/D a_n41_n33#
+ a_118_n33# w_n138_n63# pmos_5p043105913020100_3v1024x8m81_0/S_uq0 pmos_5p043105913020100_3v1024x8m81_0/S
+ pmos_5p043105913020100_3v1024x8m81
.ends

.subckt nmos_5p043105913020102_3v1024x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.353p pd=7.03u as=1.353p ps=7.03u w=3.075u l=0.28u
.ends

.subckt nmos_1p2_01_R270_3v1024x8m81 nmos_5p043105913020102_3v1024x8m81_0/D a_n14_n33#
+ nmos_5p043105913020102_3v1024x8m81_0/S VSUBS
Xnmos_5p043105913020102_3v1024x8m81_0 nmos_5p043105913020102_3v1024x8m81_0/D a_n14_n33#
+ nmos_5p043105913020102_3v1024x8m81_0/S VSUBS nmos_5p043105913020102_3v1024x8m81
.ends

.subckt xdec32_468_3v1024x8m81 LWL[6] LWL[7] RWL[18] RWL[17] RWL[15] RWL[14] RWL[13]
+ LWL[9] LWL[8] LWL[0] LWL[1] LWL[2] LWL[3] LWL[4] LWL[5] RWL[11] RWL[10] RWL[9] RWL[8]
+ RWL[7] RWL[5] RWL[1] RWL[0] LWL[18] LWL[17] LWL[16] LWL[15] LWL[14] LWL[13] LWL[12]
+ LWL[11] LWL[10] RWL[4] LWL[28] LWL[27] LWL[26] LWL[25] LWL[24] LWL[23] LWL[22] LWL[21]
+ LWL[20] LWL[19] RWL[22] RWL[26] RWL[27] RWL[30] RWL[31] LWL[31] LWL[30] LWL[29]
+ xb[3] xb[2] xb[1] xb[0] RWL[23] RWL[20] RWL[24] xa[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7219_n156#
+ RWL[21] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7483_n156# RWL[2] RWL[25] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_8012_n156#
+ xa[5] xa[4] RWL[28] RWL[12] xc RWL[3] xa[1] men xa[7] RWL[19] xa[6] RWL[16] xa[2]
+ RWL[6] RWL[29] xa[3] vdd vss
Xxdec8_3v1024x8m81_0 LWL[28] LWL[26] RWL[29] RWL[26] RWL[30] LWL[25] LWL[31] LWL[30]
+ LWL[24] LWL[27] RWL[27] xc xb[3] xa[4] xa[7] xb[3] xc xc xc xc xb[3] xa[1] xa[1]
+ RWL[24] xb[3] xc xb[1] xb[3] xa[3] xb[3] xa[0] xa[6] xa[7] RWL[25] xa[6] xb[3] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_8012_n156#
+ RWL[31] LWL[29] xc xc xb[3] xa[3] xb[2] RWL[28] xb[3] xa[5] xa[5] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7219_n156#
+ xa[2] xa[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7483_n156# men xb[0] xc xa[2]
+ xa[4] vdd vss xdec8_3v1024x8m81
Xxdec8_3v1024x8m81_1 LWL[4] LWL[2] RWL[5] RWL[2] RWL[6] LWL[1] LWL[7] LWL[6] LWL[0]
+ LWL[3] RWL[3] xc xb[0] xa[4] xa[7] xb[0] xc xc xc xc xb[0] xa[1] xa[1] RWL[0] xb[0]
+ xc xb[1] xb[0] xa[3] xb[0] xa[0] xa[6] xa[7] RWL[1] xa[6] xb[3] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_8012_n156#
+ RWL[7] LWL[5] xc xc xb[0] xa[3] xb[2] RWL[4] xb[0] xa[5] xa[5] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7219_n156#
+ xa[2] xa[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7483_n156# men xb[0] xc xa[2]
+ xa[4] vdd vss xdec8_3v1024x8m81
Xxdec8_3v1024x8m81_2 LWL[12] LWL[10] RWL[13] RWL[10] RWL[14] LWL[9] LWL[15] LWL[14]
+ LWL[8] LWL[11] RWL[11] xc xb[1] xa[4] xa[7] xb[1] xc xc xc xc xb[1] xa[1] xa[1]
+ RWL[8] xb[1] xc xb[1] xb[1] xa[3] xb[1] xa[0] xa[6] xa[7] RWL[9] xa[6] xb[3] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_8012_n156#
+ RWL[15] LWL[13] xc xc xb[1] xa[3] xb[2] RWL[12] xb[1] xa[5] xa[5] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7219_n156#
+ xa[2] xa[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7483_n156# men xb[0] xc xa[2]
+ xa[4] vdd vss xdec8_3v1024x8m81
Xxdec8_3v1024x8m81_3 LWL[20] LWL[18] RWL[21] RWL[18] RWL[22] LWL[17] LWL[23] LWL[22]
+ LWL[16] LWL[19] RWL[19] xc xb[2] xa[4] xa[7] xb[2] xc xc xc xc xb[2] xa[1] xa[1]
+ RWL[16] xb[2] xc xb[1] xb[2] xa[3] xb[2] xa[0] xa[6] xa[7] RWL[17] xa[6] xb[3] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_8012_n156#
+ RWL[23] LWL[21] xc xc xb[2] xa[3] xb[2] RWL[20] xb[2] xa[5] xa[5] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7219_n156#
+ xa[2] xa[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7483_n156# men xb[0] xc xa[2]
+ xa[4] vdd vss xdec8_3v1024x8m81
.ends

.subckt xdec64_3v1024x8m81 LWL[6] LWL[7] RWL[18] RWL[17] RWL[15] RWL[14] RWL[13] LWL[9]
+ LWL[8] LWL[0] LWL[1] LWL[2] LWL[3] LWL[4] LWL[5] RWL[11] RWL[10] RWL[9] RWL[8] RWL[7]
+ RWL[5] RWL[1] LWL[18] LWL[17] LWL[16] LWL[15] LWL[14] LWL[13] LWL[12] LWL[11] LWL[10]
+ RWL[4] LWL[28] LWL[27] LWL[26] LWL[25] LWL[24] LWL[23] LWL[22] LWL[21] LWL[20] LWL[19]
+ RWL[22] RWL[26] RWL[27] RWL[30] RWL[31] LWL[31] LWL[30] LWL[29] xa[6] xa[7] xb[3]
+ xb[2] xb[1] xb[0] RWL[23] RWL[20] xa[3] RWL[24] xa[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7219_n156#
+ RWL[21] RWL[2] RWL[25] xc xa[5] xa[4] RWL[28] RWL[12] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7748_n156#
+ RWL[3] men xa[1] RWL[19] RWL[0] xdec8_3v1024x8m81_3/xc RWL[16] xa[2] RWL[6] RWL[29]
+ vdd vss
Xxdec8_3v1024x8m81_0 LWL[28] LWL[26] RWL[29] RWL[26] RWL[30] LWL[25] LWL[31] LWL[30]
+ LWL[24] LWL[27] RWL[27] xdec8_3v1024x8m81_3/xc xb[3] xa[4] xa[7] xb[3] xdec8_3v1024x8m81_3/xc
+ xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xb[3] xa[1]
+ xa[1] RWL[24] xb[3] xdec8_3v1024x8m81_3/xc xb[1] xb[3] xa[3] xb[3] xa[0] xa[6] xa[7]
+ RWL[25] xa[6] xb[3] xc RWL[31] LWL[29] xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc
+ xb[3] xa[3] xb[2] RWL[28] xb[3] xa[5] xa[5] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7219_n156#
+ xa[2] xa[0] xdec8_3v1024x8m81_3/xc men xb[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7748_n156#
+ xa[2] xa[4] vdd vss xdec8_3v1024x8m81
Xxdec8_3v1024x8m81_1 LWL[4] LWL[2] RWL[5] RWL[2] RWL[6] LWL[1] LWL[7] LWL[6] LWL[0]
+ LWL[3] RWL[3] xdec8_3v1024x8m81_3/xc xb[0] xa[4] xa[7] xb[0] xdec8_3v1024x8m81_3/xc
+ xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xb[0] xa[1]
+ xa[1] RWL[0] xb[0] xdec8_3v1024x8m81_3/xc xb[1] xb[0] xa[3] xb[0] xa[0] xa[6] xa[7]
+ RWL[1] xa[6] xb[3] xc RWL[7] LWL[5] xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc
+ xb[0] xa[3] xb[2] RWL[4] xb[0] xa[5] xa[5] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7219_n156#
+ xa[2] xa[0] xdec8_3v1024x8m81_3/xc men xb[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7748_n156#
+ xa[2] xa[4] vdd vss xdec8_3v1024x8m81
Xxdec8_3v1024x8m81_2 LWL[12] LWL[10] RWL[13] RWL[10] RWL[14] LWL[9] LWL[15] LWL[14]
+ LWL[8] LWL[11] RWL[11] xdec8_3v1024x8m81_3/xc xb[1] xa[4] xa[7] xb[1] xdec8_3v1024x8m81_3/xc
+ xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xb[1] xa[1]
+ xa[1] RWL[8] xb[1] xdec8_3v1024x8m81_3/xc xb[1] xb[1] xa[3] xb[1] xa[0] xa[6] xa[7]
+ RWL[9] xa[6] xb[3] xc RWL[15] LWL[13] xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc
+ xb[1] xa[3] xb[2] RWL[12] xb[1] xa[5] xa[5] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7219_n156#
+ xa[2] xa[0] xdec8_3v1024x8m81_3/xc men xb[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7748_n156#
+ xa[2] xa[4] vdd vss xdec8_3v1024x8m81
Xxdec8_3v1024x8m81_3 LWL[20] LWL[18] RWL[21] RWL[18] RWL[22] LWL[17] LWL[23] LWL[22]
+ LWL[16] LWL[19] RWL[19] xdec8_3v1024x8m81_3/xc xb[2] xa[4] xa[7] xb[2] xdec8_3v1024x8m81_3/xc
+ xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc xb[2] xa[1]
+ xa[1] RWL[16] xb[2] xdec8_3v1024x8m81_3/xc xb[1] xb[2] xa[3] xb[2] xa[0] xa[6] xa[7]
+ RWL[17] xa[6] xb[3] xc RWL[23] LWL[21] xdec8_3v1024x8m81_3/xc xdec8_3v1024x8m81_3/xc
+ xb[2] xa[3] xb[2] RWL[20] xb[2] xa[5] xa[5] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7219_n156#
+ xa[2] xa[0] xdec8_3v1024x8m81_3/xc men xb[0] xdec8_3v1024x8m81_3/xdec_3v1024x8m81_7/m2_7748_n156#
+ xa[2] xa[4] vdd vss xdec8_3v1024x8m81
.ends

.subckt xdec128_3v1024x8m81 DRWL RWL[35] RWL[36] RWL[37] RWL[38] RWL[39] RWL[44] RWL[46]
+ RWL[47] RWL[48] RWL[50] RWL[51] RWL[53] RWL[54] RWL[55] RWL[56] RWL[57] RWL[58]
+ RWL[62] LWL[59] LWL[58] LWL[57] LWL[56] LWL[55] LWL[54] LWL[53] LWL[52] LWL[50]
+ LWL[45] LWL[40] LWL[38] LWL[37] LWL[36] LWL[35] LWL[34] LWL[33] DLWL LWL[19] LWL[20]
+ LWL[21] LWL[22] LWL[12] LWL[14] LWL[15] LWL[16] LWL[17] LWL[5] LWL[3] LWL[0] LWL[8]
+ LWL[9] LWL[6] LWL[29] LWL[30] RWL[32] RWL[25] RWL[6] RWL[4] RWL[2] RWL[3] RWL[5]
+ RWL[8] RWL[9] RWL[10] RWL[11] RWL[12] RWL[13] RWL[17] RWL[18] RWL[19] RWL[20] xb[0]
+ xb[1] xb[2] xb[3] xa[7] xa[6] xa[5] xa[4] xa[0] men xa[3] xa[2] xa[1] xc[0] xc[1]
+ RWL[64] RWL[65] RWL[66] RWL[69] RWL[71] RWL[72] RWL[73] RWL[74] RWL[82] RWL[84]
+ RWL[85] RWL[86] RWL[89] RWL[90] RWL[91] RWL[97] RWL[103] RWL[106] RWL[108] RWL[110]
+ RWL[111] RWL[112] RWL[113] RWL[115] RWL[116] RWL[117] RWL[118] RWL[119] RWL[123]
+ RWL[126] RWL[127] LWL[64] LWL[65] LWL[69] LWL[71] LWL[73] LWL[74] LWL[75] LWL[76]
+ LWL[77] LWL[78] LWL[79] LWL[82] LWL[84] LWL[85] LWL[89] LWL[91] LWL[92] LWL[93]
+ LWL[94] LWL[95] LWL[96] LWL[97] LWL[98] LWL[99] LWL[105] LWL[108] LWL[109] LWL[110]
+ LWL[111] LWL[112] LWL[114] LWL[115] LWL[117] LWL[118] LWL[119] RWL[93] RWL[59] RWL[92]
+ LWL[28] LWL[81] LWL[63] LWL[101] RWL[94] LWL[66] LWL[26] RWL[23] RWL[79] LWL[43]
+ RWL[75] LWL[86] LWL[100] RWL[42] LWL[27] LWL[24] LWL[120] RWL[45] RWL[76] LWL[125]
+ RWL[60] RWL[100] RWL[96] LWL[121] RWL[40] RWL[81] LWL[10] RWL[109] LWL[68] RWL[120]
+ RWL[105] LWL[61] LWL[67] RWL[99] LWL[48] RWL[101] RWL[95] LWL[88] LWL[13] LWL[102]
+ RWL[21] RWL[63] RWL[68] LWL[122] RWL[29] LWL[41] RWL[0] RWL[78] RWL[88] LWL[25]
+ RWL[102] RWL[1] RWL[98] RWL[28] LWL[1] RWL[43] RWL[122] RWL[125] LWL[87] RWL[30]
+ RWL[121] LWL[83] LWL[51] LWL[46] xdec64_468_3v1024x8m81_0/xdec8_3v1024x8m81_3/xc
+ LWL[104] RWL[26] LWL[107] RWL[67] xdec64_3v1024x8m81_0/xdec8_3v1024x8m81_3/xc LWL[124]
+ LWL[103] RWL[33] LWL[11] LWL[70] LWL[18] LWL[80] LWL[44] RWL[61] RWL[104] LWL[90]
+ RWL[24] RWL[27] LWL[39] RWL[77] RWL[114] RWL[34] LWL[4] LWL[113] RWL[124] LWL[47]
+ RWL[16] LWL[23] RWL[70] LWL[62] RWL[31] LWL[31] RWL[41] RWL[80] LWL[42] LWL[106]
+ RWL[7] RWL[52] RWL[22] LWL[7] LWL[127] RWL[49] RWL[87] LWL[116] vdd RWL[15] LWL[32]
+ LWL[2] LWL[126] LWL[123] RWL[14] RWL[83] LWL[49] LWL[72] LWL[60] RWL[107] vss
Xxdec64_468_3v1024x8m81_0 LWL[102] LWL[103] RWL[114] RWL[113] RWL[111] RWL[110] RWL[109]
+ LWL[105] LWL[104] LWL[96] LWL[97] LWL[98] LWL[99] LWL[100] LWL[101] RWL[107] RWL[106]
+ RWL[105] RWL[104] RWL[103] RWL[101] RWL[97] RWL[96] LWL[114] LWL[113] LWL[112] LWL[111]
+ LWL[110] LWL[109] LWL[108] LWL[107] LWL[106] RWL[100] LWL[124] LWL[123] LWL[122]
+ LWL[121] LWL[120] LWL[119] LWL[118] LWL[117] LWL[116] LWL[115] RWL[118] RWL[122]
+ RWL[123] RWL[126] RWL[127] LWL[127] LWL[126] LWL[125] xa[0] xa[3] xa[4] xa[5] xa[6]
+ xa[7] xb[3] xb[2] xb[1] xb[0] xc[1] xa[1] xc[0] RWL[119] RWL[116] RWL[120] RWL[117]
+ xdec64_3v1024x8m81_0/xdec8_3v1024x8m81_3/xc xa[2] RWL[98] RWL[121] RWL[124] RWL[108]
+ RWL[99] men RWL[115] xdec64_468_3v1024x8m81_0/xdec8_3v1024x8m81_3/xc RWL[112] RWL[102]
+ RWL[125] vdd vss xdec64_468_3v1024x8m81
Xnmos_5p043105913020111_3v1024x8m81_0 vss pmos_5p043105913020101_3v1024x8m81_1/D nmos_5p043105913020111_3v1024x8m81_0/S
+ vss nmos_5p043105913020111_3v1024x8m81
Xnmos_5p043105913020111_3v1024x8m81_1 vss pmos_5p043105913020101_3v1024x8m81_1/D pmos_5p043105913020101_3v1024x8m81_0/S
+ vss nmos_5p043105913020111_3v1024x8m81
Xpmos_5p043105913020101_3v1024x8m81_0 vdd pmos_5p043105913020101_3v1024x8m81_1/D vdd
+ pmos_5p043105913020101_3v1024x8m81_0/S pmos_5p043105913020101_3v1024x8m81
Xpmos_1p2_01_R90_3v1024x8m81_0 nmos_5p043105913020111_3v1024x8m81_0/S vdd pmos_5p043105913020101_3v1024x8m81_1/D
+ vdd pmos_1p2_01_R90_3v1024x8m81
Xpmos_5p043105913020101_3v1024x8m81_1 pmos_5p043105913020101_3v1024x8m81_1/D vss vdd
+ men pmos_5p043105913020101_3v1024x8m81
Xnmos_1p2_02_R90_3v1024x8m81_0 DLWL vss nmos_5p043105913020111_3v1024x8m81_0/S vss
+ nmos_1p2_02_R90_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_90 LWL[90] vss vdd LWL[91] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_91 RWL[90] vss vdd RWL[91] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_80 LWL[80] vss vdd LWL[81] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_70 LWL[70] vss vdd LWL[71] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_81 RWL[80] vss vdd RWL[81] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_92 LWL[92] vss vdd LWL[93] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_0 RWL[16] vss vdd RWL[17] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_93 RWL[92] vss vdd RWL[93] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_60 RWL[36] vss vdd RWL[37] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_71 RWL[70] vss vdd RWL[71] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_82 LWL[82] vss vdd LWL[83] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_1 RWL[14] vss vdd RWL[15] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_61 RWL[34] vss vdd RWL[35] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_50 RWL[56] vss vdd RWL[57] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_72 LWL[72] vss vdd LWL[73] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_83 RWL[82] vss vdd RWL[83] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_94 LWL[94] vss vdd LWL[95] vdd pmoscap_R270_3v1024x8m81
Xnmos_5p04310591302099_3v1024x8m81_0 vss pmos_5p043105913020101_3v1024x8m81_0/S DRWL
+ vss nmos_5p04310591302099_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_2 RWL[12] vss vdd RWL[13] vdd pmoscap_R270_3v1024x8m81
Xxdec32_3v1024x8m81_0 LWL[6] LWL[7] RWL[18] RWL[17] RWL[15] RWL[14] RWL[13] LWL[9]
+ LWL[8] LWL[0] LWL[1] LWL[2] LWL[3] LWL[4] LWL[5] RWL[11] RWL[10] RWL[9] RWL[8] RWL[7]
+ RWL[5] RWL[1] LWL[18] LWL[17] LWL[16] LWL[15] LWL[14] LWL[13] LWL[12] LWL[11] LWL[10]
+ RWL[4] LWL[28] LWL[27] LWL[26] LWL[25] LWL[24] LWL[23] LWL[22] LWL[21] LWL[20] LWL[19]
+ RWL[22] RWL[23] RWL[26] RWL[27] RWL[30] RWL[31] LWL[31] LWL[30] LWL[29] xb[3] xb[2]
+ xb[1] xb[0] RWL[20] RWL[24] xa[0] xdec64_468_3v1024x8m81_0/xdec8_3v1024x8m81_3/xc
+ RWL[21] xdec64_3v1024x8m81_0/xdec8_3v1024x8m81_3/xc RWL[2] RWL[25] xc[0] xa[5] xa[4]
+ RWL[28] RWL[12] xc[1] RWL[3] men xa[1] xa[7] RWL[19] RWL[0] xa[6] RWL[16] xa[2]
+ RWL[6] vdd RWL[29] xa[3] vss xdec32_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_95 RWL[94] vss vdd RWL[95] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_62 LWL[32] vss vdd LWL[33] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_40 LWL[46] vss vdd LWL[47] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_51 RWL[54] vss vdd RWL[55] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_73 RWL[72] vss vdd RWL[73] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_84 LWL[84] vss vdd LWL[85] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_3 RWL[10] vss vdd RWL[11] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_96 LWL[96] vss vdd LWL[97] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_30 LWL[20] vss vdd LWL[21] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_63 RWL[32] vss vdd RWL[33] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_41 LWL[44] vss vdd LWL[45] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_52 RWL[52] vss vdd RWL[53] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_74 LWL[74] vss vdd LWL[75] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_85 RWL[84] vss vdd RWL[85] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_4 RWL[8] vss vdd RWL[9] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_97 RWL[96] vss vdd RWL[97] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_20 LWL[8] vss vdd LWL[9] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_31 LWL[18] vss vdd LWL[19] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_42 LWL[42] vss vdd LWL[43] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_53 RWL[50] vss vdd RWL[51] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_64 LWL[64] vss vdd LWL[65] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_75 RWL[74] vss vdd RWL[75] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_86 LWL[86] vss vdd LWL[87] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_5 RWL[6] vss vdd RWL[7] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_98 LWL[98] vss vdd LWL[99] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_21 LWL[6] vss vdd LWL[7] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_10 RWL[28] vss vdd RWL[29] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_43 LWL[40] vss vdd LWL[41] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_54 RWL[48] vss vdd RWL[49] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_32 LWL[62] vss vdd LWL[63] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_65 RWL[64] vss vdd RWL[65] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_76 LWL[76] vss vdd LWL[77] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_87 RWL[86] vss vdd RWL[87] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_6 RWL[4] vss vdd RWL[5] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_22 LWL[4] vss vdd LWL[5] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_11 RWL[26] vss vdd RWL[27] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_44 LWL[38] vss vdd LWL[39] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_55 RWL[46] vss vdd RWL[47] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_33 LWL[60] vss vdd LWL[61] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_120 LWL[120] vss vdd LWL[121] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_99 RWL[98] vss vdd RWL[99] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_66 LWL[66] vss vdd LWL[67] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_77 RWL[76] vss vdd RWL[77] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_88 LWL[88] vss vdd LWL[89] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_7 RWL[2] vss vdd RWL[3] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_23 LWL[2] vss vdd LWL[3] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_12 RWL[24] vss vdd RWL[25] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_45 LWL[36] vss vdd LWL[37] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_56 RWL[44] vss vdd RWL[45] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_34 LWL[58] vss vdd LWL[59] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_67 RWL[66] vss vdd RWL[67] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_78 LWL[78] vss vdd LWL[79] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_89 RWL[88] vss vdd RWL[89] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_121 RWL[120] vss vdd RWL[121] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_110 LWL[110] vss vdd LWL[111] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_8 RWL[0] vss vdd RWL[1] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_L1_W2_R270_3v1024x8m81_0 DLWL vdd vss vdd vdd vdd pmoscap_L1_W2_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_122 LWL[122] vss vdd LWL[123] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_111 RWL[110] vss vdd RWL[111] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_100 LWL[100] vss vdd LWL[101] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_24 LWL[0] vss vdd LWL[1] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_13 RWL[22] vss vdd RWL[23] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_46 LWL[34] vss vdd LWL[35] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_57 RWL[42] vss vdd RWL[43] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_35 LWL[56] vss vdd LWL[57] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_68 LWL[68] vss vdd LWL[69] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_79 RWL[78] vss vdd RWL[79] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_9 RWL[30] vss vdd RWL[31] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_L1_W2_R270_3v1024x8m81_1 DRWL vdd vss vdd vdd vdd pmoscap_L1_W2_R270_3v1024x8m81
Xpmos_1p2_02_R90_3v1024x8m81_0 vdd vdd vdd nmos_5p043105913020111_3v1024x8m81_0/S
+ DLWL nmos_5p043105913020111_3v1024x8m81_0/S pmos_1p2_02_R90_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_14 RWL[20] vss vdd RWL[21] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_25 LWL[30] vss vdd LWL[31] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_58 RWL[40] vss vdd RWL[41] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_36 LWL[54] vss vdd LWL[55] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_47 RWL[62] vss vdd RWL[63] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_69 RWL[68] vss vdd RWL[69] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_123 RWL[122] vss vdd RWL[123] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_112 LWL[112] vss vdd LWL[113] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_101 RWL[100] vss vdd RWL[101] vdd pmoscap_R270_3v1024x8m81
Xpmos_1p2_02_R90_3v1024x8m81_1 vdd vdd vdd pmos_5p043105913020101_3v1024x8m81_0/S
+ DRWL pmos_5p043105913020101_3v1024x8m81_0/S pmos_1p2_02_R90_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_15 RWL[18] vss vdd RWL[19] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_26 LWL[28] vss vdd LWL[29] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_59 RWL[38] vss vdd RWL[39] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_37 LWL[52] vss vdd LWL[53] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_48 RWL[60] vss vdd RWL[61] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_124 LWL[124] vss vdd LWL[125] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_113 RWL[112] vss vdd RWL[113] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_102 LWL[102] vss vdd LWL[103] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_16 LWL[16] vss vdd LWL[17] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_27 LWL[26] vss vdd LWL[27] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_38 LWL[50] vss vdd LWL[51] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_49 RWL[58] vss vdd RWL[59] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_125 RWL[124] vss vdd RWL[125] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_114 LWL[114] vss vdd LWL[115] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_103 RWL[102] vss vdd RWL[103] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_17 LWL[14] vss vdd LWL[15] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_28 LWL[24] vss vdd LWL[25] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_39 LWL[48] vss vdd LWL[49] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_126 LWL[126] vss vdd LWL[127] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_115 RWL[114] vss vdd RWL[115] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_104 LWL[104] vss vdd LWL[105] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_18 LWL[12] vss vdd LWL[13] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_29 LWL[22] vss vdd LWL[23] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_127 RWL[126] vss vdd RWL[127] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_116 LWL[116] vss vdd LWL[117] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_105 RWL[104] vss vdd RWL[105] vdd pmoscap_R270_3v1024x8m81
Xnmos_1p2_01_R270_3v1024x8m81_0 men vdd pmos_5p043105913020101_3v1024x8m81_1/D vss
+ nmos_1p2_01_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_19 LWL[10] vss vdd LWL[11] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_117 RWL[116] vss vdd RWL[117] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_106 LWL[106] vss vdd LWL[107] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_118 LWL[118] vss vdd LWL[119] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_107 RWL[106] vss vdd RWL[107] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_119 RWL[118] vss vdd RWL[119] vdd pmoscap_R270_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_108 LWL[108] vss vdd LWL[109] vdd pmoscap_R270_3v1024x8m81
Xxdec32_468_3v1024x8m81_0 LWL[38] LWL[39] RWL[50] RWL[49] RWL[47] RWL[46] RWL[45]
+ LWL[41] LWL[40] LWL[32] LWL[33] LWL[34] LWL[35] LWL[36] LWL[37] RWL[43] RWL[42]
+ RWL[41] RWL[40] RWL[39] RWL[37] RWL[33] RWL[32] LWL[50] LWL[49] LWL[48] LWL[47]
+ LWL[46] LWL[45] LWL[44] LWL[43] LWL[42] RWL[36] LWL[60] LWL[59] LWL[58] LWL[57]
+ LWL[56] LWL[55] LWL[54] LWL[53] LWL[52] LWL[51] RWL[54] RWL[58] RWL[59] RWL[62]
+ RWL[63] LWL[63] LWL[62] LWL[61] xb[3] xb[2] xb[1] xb[0] RWL[55] RWL[52] RWL[56]
+ xa[0] xdec64_468_3v1024x8m81_0/xdec8_3v1024x8m81_3/xc RWL[53] xdec64_3v1024x8m81_0/xdec8_3v1024x8m81_3/xc
+ RWL[34] RWL[57] xc[0] xa[5] xa[4] RWL[60] RWL[44] xc[1] RWL[35] xa[1] men xa[7]
+ RWL[51] xa[6] RWL[48] xa[2] RWL[38] RWL[61] xa[3] vdd vss xdec32_468_3v1024x8m81
Xpmoscap_R270_3v1024x8m81_109 RWL[108] vss vdd RWL[109] vdd pmoscap_R270_3v1024x8m81
Xxdec64_3v1024x8m81_0 LWL[70] LWL[71] RWL[82] RWL[81] RWL[79] RWL[78] RWL[77] LWL[73]
+ LWL[72] LWL[64] LWL[65] LWL[66] LWL[67] LWL[68] LWL[69] RWL[75] RWL[74] RWL[73]
+ RWL[72] RWL[71] RWL[69] RWL[65] LWL[82] LWL[81] LWL[80] LWL[79] LWL[78] LWL[77]
+ LWL[76] LWL[75] LWL[74] RWL[68] LWL[92] LWL[91] LWL[90] LWL[89] LWL[88] LWL[87]
+ LWL[86] LWL[85] LWL[84] LWL[83] RWL[86] RWL[90] RWL[91] RWL[94] RWL[95] LWL[95]
+ LWL[94] LWL[93] xa[6] xa[7] xb[3] xb[2] xb[1] xb[0] RWL[87] RWL[84] xa[3] RWL[88]
+ xa[0] xdec64_468_3v1024x8m81_0/xdec8_3v1024x8m81_3/xc RWL[85] RWL[66] RWL[89] xc[0]
+ xa[5] xa[4] RWL[92] RWL[76] xc[1] RWL[67] men xa[1] RWL[83] RWL[64] xdec64_3v1024x8m81_0/xdec8_3v1024x8m81_3/xc
+ RWL[80] xa[2] RWL[70] RWL[93] vdd vss xdec64_3v1024x8m81
.ends

.subckt gf180mcu_ocd_ip_sram__sram1024x8m8wm1 A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1]
+ A[0] CEN CLK D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] GWEN Q[7] Q[6] Q[5] Q[4] Q[3]
+ Q[2] Q[1] Q[0] VDD VSS WEN[7] WEN[6] WEN[5] WEN[4] WEN[3] WEN[2] WEN[1] WEN[0] A[9]
Xrcol4_1024_3v1024x8m81_0 xdec128_3v1024x8m81_0/RWL[33] rcol4_1024_3v1024x8m81_0/WL[33]
+ xdec128_3v1024x8m81_0/RWL[35] rcol4_1024_3v1024x8m81_0/WL[35] xdec128_3v1024x8m81_0/RWL[37]
+ VSS xdec128_3v1024x8m81_0/RWL[50] xdec128_3v1024x8m81_0/RWL[52] xdec128_3v1024x8m81_0/RWL[54]
+ xdec128_3v1024x8m81_0/RWL[56] rcol4_1024_3v1024x8m81_0/WL[56] xdec128_3v1024x8m81_0/RWL[63]
+ xdec128_3v1024x8m81_0/RWL[53] xdec128_3v1024x8m81_0/RWL[30] xdec128_3v1024x8m81_0/RWL[26]
+ xdec128_3v1024x8m81_0/RWL[25] rcol4_1024_3v1024x8m81_0/WL[20] xdec128_3v1024x8m81_0/RWL[28]
+ xdec128_3v1024x8m81_0/RWL[31] VSS VSS xdec128_3v1024x8m81_0/RWL[16] rcol4_1024_3v1024x8m81_0/WL[38]
+ rcol4_1024_3v1024x8m81_0/WL[45] VSS xdec128_3v1024x8m81_0/RWL[42] VSS rcol4_1024_3v1024x8m81_0/WL[31]
+ VSS VSS xdec128_3v1024x8m81_0/RWL[18] xdec128_3v1024x8m81_0/RWL[27] xdec128_3v1024x8m81_0/RWL[20]
+ rcol4_1024_3v1024x8m81_0/WL[58] rcol4_1024_3v1024x8m81_0/WL[60] rcol4_1024_3v1024x8m81_0/WL[62]
+ xdec128_3v1024x8m81_0/RWL[55] xdec128_3v1024x8m81_0/RWL[49] xdec128_3v1024x8m81_0/RWL[57]
+ VSS rcol4_1024_3v1024x8m81_0/WL[8] xdec128_3v1024x8m81_0/RWL[5] VSS rcol4_1024_3v1024x8m81_0/WL[13]
+ rcol4_1024_3v1024x8m81_0/WL[6] rcol4_1024_3v1024x8m81_0/tblhl rcol4_1024_3v1024x8m81_0/GWE
+ xdec128_3v1024x8m81_0/RWL[11] D[7] Q[5] Q[6] Q[7] D[5] D[6] Q[4] rcol4_1024_3v1024x8m81_0/pcb[6]
+ rcol4_1024_3v1024x8m81_0/pcb[7] WEN[7] WEN[4] rcol4_1024_3v1024x8m81_0/pcb[5] WEN[6]
+ WEN[5] D[4] xdec128_3v1024x8m81_0/RWL[41] xdec128_3v1024x8m81_0/RWL[69] xdec128_3v1024x8m81_0/RWL[40]
+ xdec128_3v1024x8m81_0/RWL[99] xdec128_3v1024x8m81_0/RWL[68] xdec128_3v1024x8m81_0/RWL[14]
+ xdec128_3v1024x8m81_0/RWL[113] rcol4_1024_3v1024x8m81_0/pcb[4] xdec128_3v1024x8m81_0/RWL[94]
+ xdec128_3v1024x8m81_0/RWL[13] xdec128_3v1024x8m81_0/RWL[122] xdec128_3v1024x8m81_0/RWL[79]
+ xdec128_3v1024x8m81_0/RWL[107] xdec128_3v1024x8m81_0/RWL[78] xdec128_3v1024x8m81_0/RWL[106]
+ xdec128_3v1024x8m81_0/RWL[121] xdec128_3v1024x8m81_0/RWL[34] xdec128_3v1024x8m81_0/RWL[17]
+ xdec128_3v1024x8m81_0/RWL[0] xdec128_3v1024x8m81_0/RWL[71] xdec128_3v1024x8m81_0/RWL[115]
+ xdec128_3v1024x8m81_0/RWL[70] xdec128_3v1024x8m81_0/RWL[100] xdec128_3v1024x8m81_0/RWL[83]
+ xdec128_3v1024x8m81_0/RWL[15] xdec128_3v1024x8m81_0/RWL[124] xdec128_3v1024x8m81_0/RWL[21]
+ xdec128_3v1024x8m81_0/RWL[81] xdec128_3v1024x8m81_0/RWL[109] xdec128_3v1024x8m81_0/RWL[80]
+ xdec128_3v1024x8m81_0/RWL[108] xdec128_3v1024x8m81_0/RWL[8] xdec128_3v1024x8m81_0/RWL[65]
+ xdec128_3v1024x8m81_0/RWL[19] xdec128_3v1024x8m81_0/RWL[93] xdec128_3v1024x8m81_0/RWL[74]
+ xdec128_3v1024x8m81_0/RWL[102] xdec128_3v1024x8m81_0/RWL[7] xdec128_3v1024x8m81_0/RWL[59]
+ xdec128_3v1024x8m81_0/RWL[87] xdec128_3v1024x8m81_0/RWL[6] xdec128_3v1024x8m81_0/RWL[58]
+ xdec128_3v1024x8m81_0/RWL[101] xdec128_3v1024x8m81_0/RWL[86] xdec128_3v1024x8m81_0/RWL[44]
+ VSS xdec128_3v1024x8m81_0/RWL[72] xdec128_3v1024x8m81_0/RWL[1] xdec128_3v1024x8m81_0/RWL[116]
+ xdec128_3v1024x8m81_0/RWL[43] xdec128_3v1024x8m81_0/RWL[29] xdec128_3v1024x8m81_0/RWL[85]
+ xdec128_3v1024x8m81_0/RWL[112] xdec128_3v1024x8m81_0/RWL[97] rcol4_1024_3v1024x8m81_0/pcb[4]
+ xdec128_3v1024x8m81_0/RWL[51] xdec128_3v1024x8m81_0/RWL[36] xdec128_3v1024x8m81_0/RWL[125]
+ xdec128_3v1024x8m81_0/RWL[22] xdec128_3v1024x8m81_0/RWL[96] xdec128_3v1024x8m81_0/RWL[111]
+ xdec128_3v1024x8m81_0/RWL[66] xdec128_3v1024x8m81_0/RWL[82] xdec128_3v1024x8m81_0/RWL[110]
+ xdec128_3v1024x8m81_0/RWL[10] xdec128_3v1024x8m81_0/DRWL xdec128_3v1024x8m81_0/RWL[95]
+ xdec128_3v1024x8m81_0/RWL[123] xdec128_3v1024x8m81_0/RWL[104] xdec128_3v1024x8m81_0/RWL[9]
+ xdec128_3v1024x8m81_0/RWL[61] xdec128_3v1024x8m81_0/RWL[46] xdec128_3v1024x8m81_0/RWL[89]
+ xdec128_3v1024x8m81_0/RWL[32] xdec128_3v1024x8m81_0/RWL[117] xdec128_3v1024x8m81_0/RWL[60]
+ xdec128_3v1024x8m81_0/RWL[88] control_3v1024x8_3v1024x8m81_0/RYS[0] xdec128_3v1024x8m81_0/RWL[45]
+ VDD xdec128_3v1024x8m81_0/RWL[73] xdec128_3v1024x8m81_0/RWL[2] control_3v1024x8_3v1024x8m81_0/RYS[1]
+ VDD xdec128_3v1024x8m81_0/RWL[114] xdec128_3v1024x8m81_0/RWL[84] control_3v1024x8_3v1024x8m81_0/RYS[2]
+ xdec128_3v1024x8m81_0/RWL[39] VDD xdec128_3v1024x8m81_0/RWL[67] xdec128_3v1024x8m81_0/RWL[38]
+ xdec128_3v1024x8m81_0/RWL[127] control_3v1024x8_3v1024x8m81_0/RYS[3] xdec128_3v1024x8m81_0/RWL[24]
+ xdec128_3v1024x8m81_0/RWL[98] xdec128_3v1024x8m81_0/RWL[126] xdec128_3v1024x8m81_0/RWL[23]
+ control_3v1024x8_3v1024x8m81_0/RYS[4] xdec128_3v1024x8m81_0/men xdec128_3v1024x8m81_0/RWL[12]
+ xdec128_3v1024x8m81_0/RWL[64] control_3v1024x8_3v1024x8m81_0/RYS[5] xdec128_3v1024x8m81_0/RWL[92]
+ VDD xdec128_3v1024x8m81_0/RWL[120] VDD control_3v1024x8_3v1024x8m81_0/RYS[6] xdec128_3v1024x8m81_0/RWL[77]
+ xdec128_3v1024x8m81_0/RWL[105] xdec128_3v1024x8m81_0/RWL[48] xdec128_3v1024x8m81_0/RWL[91]
+ xdec128_3v1024x8m81_0/RWL[76] control_3v1024x8_3v1024x8m81_0/RYS[7] xdec128_3v1024x8m81_0/RWL[119]
+ xdec128_3v1024x8m81_0/RWL[62] xdec128_3v1024x8m81_0/RWL[90] VDD control_3v1024x8_3v1024x8m81_0/IGWEN
+ xdec128_3v1024x8m81_0/RWL[118] xdec128_3v1024x8m81_0/RWL[47] xdec128_3v1024x8m81_0/RWL[75]
+ xdec128_3v1024x8m81_0/RWL[4] VDD xdec128_3v1024x8m81_0/RWL[103] VDD xdec128_3v1024x8m81_0/RWL[3]
+ VSS rcol4_1024_3v1024x8m81
Xlcol4_1024_3v1024x8m81_0 xdec128_3v1024x8m81_0/LWL[33] lcol4_1024_3v1024x8m81_0/WL[33]
+ xdec128_3v1024x8m81_0/LWL[35] lcol4_1024_3v1024x8m81_0/WL[38] VSS VSS xdec128_3v1024x8m81_0/LWL[37]
+ VSS VSS lcol4_1024_3v1024x8m81_0/WL[43] lcol4_1024_3v1024x8m81_0/WL[45] xdec128_3v1024x8m81_0/LWL[50]
+ xdec128_3v1024x8m81_0/LWL[51] xdec128_3v1024x8m81_0/LWL[52] xdec128_3v1024x8m81_0/LWL[53]
+ xdec128_3v1024x8m81_0/LWL[54] xdec128_3v1024x8m81_0/LWL[55] xdec128_3v1024x8m81_0/LWL[56]
+ xdec128_3v1024x8m81_0/LWL[57] lcol4_1024_3v1024x8m81_0/WL[56] lcol4_1024_3v1024x8m81_0/WL[58]
+ VSS lcol4_1024_3v1024x8m81_0/WL[63] lcol4_1024_3v1024x8m81_0/WL[20] xdec128_3v1024x8m81_0/LWL[20]
+ lcol4_1024_3v1024x8m81_0/WL[18] xdec128_3v1024x8m81_0/LWL[18] VSS xdec128_3v1024x8m81_0/LWL[16]
+ VSS lcol4_1024_3v1024x8m81_0/WL[13] VSS VSS xdec128_3v1024x8m81_0/LWL[9] lcol4_1024_3v1024x8m81_0/WL[8]
+ lcol4_1024_3v1024x8m81_0/WL[6] lcol4_1024_3v1024x8m81_0/WL[31] xdec128_3v1024x8m81_0/LWL[31]
+ xdec128_3v1024x8m81_0/LWL[30] D[1] D[3] D[2] Q[1] Q[2] Q[3] lcol4_1024_3v1024x8m81_0/pcb[2]
+ lcol4_1024_3v1024x8m81_0/pcb[3] lcol4_1024_3v1024x8m81_0/pcb[0] lcol4_1024_3v1024x8m81_0/pcb[1]
+ WEN[0] WEN[1] WEN[2] Q[0] D[0] xdec128_3v1024x8m81_0/LWL[76] xdec128_3v1024x8m81_0/LWL[14]
+ xdec128_3v1024x8m81_0/LWL[113] xdec128_3v1024x8m81_0/LWL[86] xdec128_3v1024x8m81_0/LWL[123]
+ xdec128_3v1024x8m81_0/LWL[15] xdec128_3v1024x8m81_0/LWL[96] xdec128_3v1024x8m81_0/LWL[32]
+ xdec128_3v1024x8m81_0/LWL[69] xdec128_3v1024x8m81_0/LWL[102] xdec128_3v1024x8m81_0/LWL[79]
+ xdec128_3v1024x8m81_0/LWL[17] xdec128_3v1024x8m81_0/LWL[34] xdec128_3v1024x8m81_0/LWL[112]
+ xdec128_3v1024x8m81_0/LWL[89] xdec128_3v1024x8m81_0/LWL[122] xdec128_3v1024x8m81_0/LWL[99]
+ xdec128_3v1024x8m81_0/LWL[19] xdec128_3v1024x8m81_0/LWL[68] xdec128_3v1024x8m81_0/LWL[36]
+ VDD xdec128_3v1024x8m81_0/LWL[105] xdec128_3v1024x8m81_0/LWL[78] xdec128_3v1024x8m81_0/LWL[115]
+ xdec128_3v1024x8m81_0/LWL[88] xdec128_3v1024x8m81_0/LWL[38] xdec128_3v1024x8m81_0/LWL[125]
+ xdec128_3v1024x8m81_0/LWL[98] xdec128_3v1024x8m81_0/LWL[39] xdec128_3v1024x8m81_0/LWL[104]
+ xdec128_3v1024x8m81_0/LWL[114] xdec128_3v1024x8m81_0/LWL[58] xdec128_3v1024x8m81_0/LWL[124]
+ xdec128_3v1024x8m81_0/LWL[59] xdec128_3v1024x8m81_0/LWL[107] xdec128_3v1024x8m81_0/LWL[71]
+ xdec128_3v1024x8m81_0/LWL[117] xdec128_3v1024x8m81_0/LWL[81] xdec128_3v1024x8m81_0/LWL[91]
+ control_3v1024x8_3v1024x8m81_0/IGWEN xdec128_3v1024x8m81_0/LWL[106] xdec128_3v1024x8m81_0/LWL[70]
+ xdec128_3v1024x8m81_0/LWL[116] xdec128_3v1024x8m81_0/LWL[21] xdec128_3v1024x8m81_0/LWL[80]
+ xdec128_3v1024x8m81_0/LWL[126] xdec128_3v1024x8m81_0/LWL[90] xdec128_3v1024x8m81_0/LWL[22]
+ control_3v1024x8_3v1024x8m81_0/LYS[0] xdec128_3v1024x8m81_0/LWL[23] xdec128_3v1024x8m81_0/LWL[40]
+ xdec128_3v1024x8m81_0/LWL[109] xdec128_3v1024x8m81_0/LWL[73] control_3v1024x8_3v1024x8m81_0/LYS[1]
+ xdec128_3v1024x8m81_0/LWL[24] xdec128_3v1024x8m81_0/LWL[119] xdec128_3v1024x8m81_0/LWL[41]
+ xdec128_3v1024x8m81_0/LWL[83] control_3v1024x8_3v1024x8m81_0/LYS[2] xdec128_3v1024x8m81_0/LWL[25]
+ xdec128_3v1024x8m81_0/LWL[93] xdec128_3v1024x8m81_0/LWL[42] control_3v1024x8_3v1024x8m81_0/LYS[3]
+ xdec128_3v1024x8m81_0/LWL[26] xdec128_3v1024x8m81_0/LWL[43] xdec128_3v1024x8m81_0/LWL[60]
+ xdec128_3v1024x8m81_0/LWL[108] xdec128_3v1024x8m81_0/LWL[72] control_3v1024x8_3v1024x8m81_0/LYS[4]
+ xdec128_3v1024x8m81_0/LWL[27] xdec128_3v1024x8m81_0/LWL[44] xdec128_3v1024x8m81_0/LWL[118]
+ xdec128_3v1024x8m81_0/LWL[61] xdec128_3v1024x8m81_0/LWL[82] control_3v1024x8_3v1024x8m81_0/LYS[5]
+ xdec128_3v1024x8m81_0/LWL[28] xdec128_3v1024x8m81_0/LWL[45] xdec128_3v1024x8m81_0/LWL[62]
+ xdec128_3v1024x8m81_0/LWL[92] control_3v1024x8_3v1024x8m81_0/LYS[6] xdec128_3v1024x8m81_0/LWL[29]
+ xdec128_3v1024x8m81_0/LWL[46] xdec128_3v1024x8m81_0/LWL[65] control_3v1024x8_3v1024x8m81_0/LYS[7]
+ xdec128_3v1024x8m81_0/LWL[75] xdec128_3v1024x8m81_0/LWL[47] xdec128_3v1024x8m81_0/LWL[85]
+ VDD xdec128_3v1024x8m81_0/LWL[127] xdec128_3v1024x8m81_0/LWL[48] xdec128_3v1024x8m81_0/LWL[0]
+ xdec128_3v1024x8m81_0/LWL[95] VDD xdec128_3v1024x8m81_0/LWL[49] xdec128_3v1024x8m81_0/LWL[64]
+ xdec128_3v1024x8m81_0/LWL[1] xdec128_3v1024x8m81_0/LWL[101] xdec128_3v1024x8m81_0/LWL[74]
+ xdec128_3v1024x8m81_0/LWL[2] xdec128_3v1024x8m81_0/LWL[111] VDD xdec128_3v1024x8m81_0/LWL[84]
+ xdec128_3v1024x8m81_0/LWL[3] xdec128_3v1024x8m81_0/LWL[121] VDD xdec128_3v1024x8m81_0/LWL[94]
+ xdec128_3v1024x8m81_0/LWL[4] xdec128_3v1024x8m81_0/LWL[67] xdec128_3v1024x8m81_0/LWL[63]
+ xdec128_3v1024x8m81_0/LWL[100] xdec128_3v1024x8m81_0/LWL[10] xdec128_3v1024x8m81_0/LWL[77]
+ xdec128_3v1024x8m81_0/LWL[5] xdec128_3v1024x8m81_0/LWL[110] xdec128_3v1024x8m81_0/LWL[11]
+ xdec128_3v1024x8m81_0/LWL[87] VDD xdec128_3v1024x8m81_0/LWL[6] xdec128_3v1024x8m81_0/LWL[120]
+ WEN[3] xdec128_3v1024x8m81_0/LWL[97] xdec128_3v1024x8m81_0/LWL[12] xdec128_3v1024x8m81_0/LWL[7]
+ VDD rcol4_1024_3v1024x8m81_0/GWE xdec128_3v1024x8m81_0/LWL[66] xdec128_3v1024x8m81_0/men
+ VDD xdec128_3v1024x8m81_0/LWL[13] VDD xdec128_3v1024x8m81_0/LWL[103] xdec128_3v1024x8m81_0/LWL[8]
+ VSS lcol4_1024_3v1024x8m81
Xcontrol_3v1024x8_3v1024x8m81_0 control_3v1024x8_3v1024x8m81_0/RYS[7] control_3v1024x8_3v1024x8m81_0/RYS[6]
+ control_3v1024x8_3v1024x8m81_0/RYS[5] control_3v1024x8_3v1024x8m81_0/RYS[4] control_3v1024x8_3v1024x8m81_0/RYS[3]
+ control_3v1024x8_3v1024x8m81_0/RYS[2] control_3v1024x8_3v1024x8m81_0/RYS[1] control_3v1024x8_3v1024x8m81_0/RYS[0]
+ control_3v1024x8_3v1024x8m81_0/LYS[0] control_3v1024x8_3v1024x8m81_0/LYS[1] control_3v1024x8_3v1024x8m81_0/LYS[2]
+ control_3v1024x8_3v1024x8m81_0/LYS[3] control_3v1024x8_3v1024x8m81_0/LYS[6] control_3v1024x8_3v1024x8m81_0/LYS[5]
+ control_3v1024x8_3v1024x8m81_0/LYS[4] control_3v1024x8_3v1024x8m81_0/LYS[7] rcol4_1024_3v1024x8m81_0/tblhl
+ control_3v1024x8_3v1024x8m81_0/IGWEN xdec128_3v1024x8m81_0/xb[3] xdec128_3v1024x8m81_0/xb[2]
+ xdec128_3v1024x8m81_0/xb[0] xdec128_3v1024x8m81_0/xa[7] xdec128_3v1024x8m81_0/xa[6]
+ xdec128_3v1024x8m81_0/xa[5] xdec128_3v1024x8m81_0/xa[4] xdec128_3v1024x8m81_0/xa[2]
+ A[0] xdec128_3v1024x8m81_0/xb[1] control_3v1024x8_3v1024x8m81_0/xc[3] control_3v1024x8_3v1024x8m81_0/xc[2]
+ xdec128_3v1024x8m81_0/xa[1] A[9] A[7] CLK A[2] A[1] A[6] A[3] A[4] A[5] A[8] GWEN
+ control_3v1024x8_3v1024x8m81_0/VDD_uq0 VDD VDD VSS VDD xdec128_3v1024x8m81_0/xa[0]
+ xdec128_3v1024x8m81_0/xa[3] xdec128_3v1024x8m81_0/men CEN VDD xdec128_3v1024x8m81_0/xc[1]
+ VDD xdec128_3v1024x8m81_0/xc[0] rcol4_1024_3v1024x8m81_0/GWE VDD VDD VSS control_3v1024x8_3v1024x8m81
Xxdec128_3v1024x8m81_0 xdec128_3v1024x8m81_0/DRWL xdec128_3v1024x8m81_0/RWL[35] xdec128_3v1024x8m81_0/RWL[36]
+ xdec128_3v1024x8m81_0/RWL[37] xdec128_3v1024x8m81_0/RWL[38] xdec128_3v1024x8m81_0/RWL[39]
+ xdec128_3v1024x8m81_0/RWL[44] xdec128_3v1024x8m81_0/RWL[46] xdec128_3v1024x8m81_0/RWL[47]
+ xdec128_3v1024x8m81_0/RWL[48] xdec128_3v1024x8m81_0/RWL[50] xdec128_3v1024x8m81_0/RWL[51]
+ xdec128_3v1024x8m81_0/RWL[53] xdec128_3v1024x8m81_0/RWL[54] xdec128_3v1024x8m81_0/RWL[55]
+ xdec128_3v1024x8m81_0/RWL[56] xdec128_3v1024x8m81_0/RWL[57] xdec128_3v1024x8m81_0/RWL[58]
+ xdec128_3v1024x8m81_0/RWL[62] xdec128_3v1024x8m81_0/LWL[59] xdec128_3v1024x8m81_0/LWL[58]
+ xdec128_3v1024x8m81_0/LWL[57] xdec128_3v1024x8m81_0/LWL[56] xdec128_3v1024x8m81_0/LWL[55]
+ xdec128_3v1024x8m81_0/LWL[54] xdec128_3v1024x8m81_0/LWL[53] xdec128_3v1024x8m81_0/LWL[52]
+ xdec128_3v1024x8m81_0/LWL[50] xdec128_3v1024x8m81_0/LWL[45] xdec128_3v1024x8m81_0/LWL[40]
+ xdec128_3v1024x8m81_0/LWL[38] xdec128_3v1024x8m81_0/LWL[37] xdec128_3v1024x8m81_0/LWL[36]
+ xdec128_3v1024x8m81_0/LWL[35] xdec128_3v1024x8m81_0/LWL[34] xdec128_3v1024x8m81_0/LWL[33]
+ xdec128_3v1024x8m81_0/DLWL xdec128_3v1024x8m81_0/LWL[19] xdec128_3v1024x8m81_0/LWL[20]
+ xdec128_3v1024x8m81_0/LWL[21] xdec128_3v1024x8m81_0/LWL[22] xdec128_3v1024x8m81_0/LWL[12]
+ xdec128_3v1024x8m81_0/LWL[14] xdec128_3v1024x8m81_0/LWL[15] xdec128_3v1024x8m81_0/LWL[16]
+ xdec128_3v1024x8m81_0/LWL[17] xdec128_3v1024x8m81_0/LWL[5] xdec128_3v1024x8m81_0/LWL[3]
+ xdec128_3v1024x8m81_0/LWL[0] xdec128_3v1024x8m81_0/LWL[8] xdec128_3v1024x8m81_0/LWL[9]
+ xdec128_3v1024x8m81_0/LWL[6] xdec128_3v1024x8m81_0/LWL[29] xdec128_3v1024x8m81_0/LWL[30]
+ xdec128_3v1024x8m81_0/RWL[32] xdec128_3v1024x8m81_0/RWL[25] xdec128_3v1024x8m81_0/RWL[6]
+ xdec128_3v1024x8m81_0/RWL[4] xdec128_3v1024x8m81_0/RWL[2] xdec128_3v1024x8m81_0/RWL[3]
+ xdec128_3v1024x8m81_0/RWL[5] xdec128_3v1024x8m81_0/RWL[8] xdec128_3v1024x8m81_0/RWL[9]
+ xdec128_3v1024x8m81_0/RWL[10] xdec128_3v1024x8m81_0/RWL[11] xdec128_3v1024x8m81_0/RWL[12]
+ xdec128_3v1024x8m81_0/RWL[13] xdec128_3v1024x8m81_0/RWL[17] xdec128_3v1024x8m81_0/RWL[18]
+ xdec128_3v1024x8m81_0/RWL[19] xdec128_3v1024x8m81_0/RWL[20] xdec128_3v1024x8m81_0/xb[0]
+ xdec128_3v1024x8m81_0/xb[1] xdec128_3v1024x8m81_0/xb[2] xdec128_3v1024x8m81_0/xb[3]
+ xdec128_3v1024x8m81_0/xa[7] xdec128_3v1024x8m81_0/xa[6] xdec128_3v1024x8m81_0/xa[5]
+ xdec128_3v1024x8m81_0/xa[4] xdec128_3v1024x8m81_0/xa[0] xdec128_3v1024x8m81_0/men
+ xdec128_3v1024x8m81_0/xa[3] xdec128_3v1024x8m81_0/xa[2] xdec128_3v1024x8m81_0/xa[1]
+ xdec128_3v1024x8m81_0/xc[0] xdec128_3v1024x8m81_0/xc[1] xdec128_3v1024x8m81_0/RWL[64]
+ xdec128_3v1024x8m81_0/RWL[65] xdec128_3v1024x8m81_0/RWL[66] xdec128_3v1024x8m81_0/RWL[69]
+ xdec128_3v1024x8m81_0/RWL[71] xdec128_3v1024x8m81_0/RWL[72] xdec128_3v1024x8m81_0/RWL[73]
+ xdec128_3v1024x8m81_0/RWL[74] xdec128_3v1024x8m81_0/RWL[82] xdec128_3v1024x8m81_0/RWL[84]
+ xdec128_3v1024x8m81_0/RWL[85] xdec128_3v1024x8m81_0/RWL[86] xdec128_3v1024x8m81_0/RWL[89]
+ xdec128_3v1024x8m81_0/RWL[90] xdec128_3v1024x8m81_0/RWL[91] xdec128_3v1024x8m81_0/RWL[97]
+ xdec128_3v1024x8m81_0/RWL[103] xdec128_3v1024x8m81_0/RWL[106] xdec128_3v1024x8m81_0/RWL[108]
+ xdec128_3v1024x8m81_0/RWL[110] xdec128_3v1024x8m81_0/RWL[111] xdec128_3v1024x8m81_0/RWL[112]
+ xdec128_3v1024x8m81_0/RWL[113] xdec128_3v1024x8m81_0/RWL[115] xdec128_3v1024x8m81_0/RWL[116]
+ xdec128_3v1024x8m81_0/RWL[117] xdec128_3v1024x8m81_0/RWL[118] xdec128_3v1024x8m81_0/RWL[119]
+ xdec128_3v1024x8m81_0/RWL[123] xdec128_3v1024x8m81_0/RWL[126] xdec128_3v1024x8m81_0/RWL[127]
+ xdec128_3v1024x8m81_0/LWL[64] xdec128_3v1024x8m81_0/LWL[65] xdec128_3v1024x8m81_0/LWL[69]
+ xdec128_3v1024x8m81_0/LWL[71] xdec128_3v1024x8m81_0/LWL[73] xdec128_3v1024x8m81_0/LWL[74]
+ xdec128_3v1024x8m81_0/LWL[75] xdec128_3v1024x8m81_0/LWL[76] xdec128_3v1024x8m81_0/LWL[77]
+ xdec128_3v1024x8m81_0/LWL[78] xdec128_3v1024x8m81_0/LWL[79] xdec128_3v1024x8m81_0/LWL[82]
+ xdec128_3v1024x8m81_0/LWL[84] xdec128_3v1024x8m81_0/LWL[85] xdec128_3v1024x8m81_0/LWL[89]
+ xdec128_3v1024x8m81_0/LWL[91] xdec128_3v1024x8m81_0/LWL[92] xdec128_3v1024x8m81_0/LWL[93]
+ xdec128_3v1024x8m81_0/LWL[94] xdec128_3v1024x8m81_0/LWL[95] xdec128_3v1024x8m81_0/LWL[96]
+ xdec128_3v1024x8m81_0/LWL[97] xdec128_3v1024x8m81_0/LWL[98] xdec128_3v1024x8m81_0/LWL[99]
+ xdec128_3v1024x8m81_0/LWL[105] xdec128_3v1024x8m81_0/LWL[108] xdec128_3v1024x8m81_0/LWL[109]
+ xdec128_3v1024x8m81_0/LWL[110] xdec128_3v1024x8m81_0/LWL[111] xdec128_3v1024x8m81_0/LWL[112]
+ xdec128_3v1024x8m81_0/LWL[114] xdec128_3v1024x8m81_0/LWL[115] xdec128_3v1024x8m81_0/LWL[117]
+ xdec128_3v1024x8m81_0/LWL[118] xdec128_3v1024x8m81_0/LWL[119] xdec128_3v1024x8m81_0/RWL[93]
+ xdec128_3v1024x8m81_0/RWL[59] xdec128_3v1024x8m81_0/RWL[92] xdec128_3v1024x8m81_0/LWL[28]
+ xdec128_3v1024x8m81_0/LWL[81] xdec128_3v1024x8m81_0/LWL[63] xdec128_3v1024x8m81_0/LWL[101]
+ xdec128_3v1024x8m81_0/RWL[94] xdec128_3v1024x8m81_0/LWL[66] xdec128_3v1024x8m81_0/LWL[26]
+ xdec128_3v1024x8m81_0/RWL[23] xdec128_3v1024x8m81_0/RWL[79] xdec128_3v1024x8m81_0/LWL[43]
+ xdec128_3v1024x8m81_0/RWL[75] xdec128_3v1024x8m81_0/LWL[86] xdec128_3v1024x8m81_0/LWL[100]
+ xdec128_3v1024x8m81_0/RWL[42] xdec128_3v1024x8m81_0/LWL[27] xdec128_3v1024x8m81_0/LWL[24]
+ xdec128_3v1024x8m81_0/LWL[120] xdec128_3v1024x8m81_0/RWL[45] xdec128_3v1024x8m81_0/RWL[76]
+ xdec128_3v1024x8m81_0/LWL[125] xdec128_3v1024x8m81_0/RWL[60] xdec128_3v1024x8m81_0/RWL[100]
+ xdec128_3v1024x8m81_0/RWL[96] xdec128_3v1024x8m81_0/LWL[121] xdec128_3v1024x8m81_0/RWL[40]
+ xdec128_3v1024x8m81_0/RWL[81] xdec128_3v1024x8m81_0/LWL[10] xdec128_3v1024x8m81_0/RWL[109]
+ xdec128_3v1024x8m81_0/LWL[68] xdec128_3v1024x8m81_0/RWL[120] xdec128_3v1024x8m81_0/RWL[105]
+ xdec128_3v1024x8m81_0/LWL[61] xdec128_3v1024x8m81_0/LWL[67] xdec128_3v1024x8m81_0/RWL[99]
+ xdec128_3v1024x8m81_0/LWL[48] xdec128_3v1024x8m81_0/RWL[101] xdec128_3v1024x8m81_0/RWL[95]
+ xdec128_3v1024x8m81_0/LWL[88] xdec128_3v1024x8m81_0/LWL[13] xdec128_3v1024x8m81_0/LWL[102]
+ xdec128_3v1024x8m81_0/RWL[21] xdec128_3v1024x8m81_0/RWL[63] xdec128_3v1024x8m81_0/RWL[68]
+ xdec128_3v1024x8m81_0/LWL[122] xdec128_3v1024x8m81_0/RWL[29] xdec128_3v1024x8m81_0/LWL[41]
+ xdec128_3v1024x8m81_0/RWL[0] xdec128_3v1024x8m81_0/RWL[78] xdec128_3v1024x8m81_0/RWL[88]
+ xdec128_3v1024x8m81_0/LWL[25] xdec128_3v1024x8m81_0/RWL[102] xdec128_3v1024x8m81_0/RWL[1]
+ xdec128_3v1024x8m81_0/RWL[98] xdec128_3v1024x8m81_0/RWL[28] xdec128_3v1024x8m81_0/LWL[1]
+ xdec128_3v1024x8m81_0/RWL[43] xdec128_3v1024x8m81_0/RWL[122] xdec128_3v1024x8m81_0/RWL[125]
+ xdec128_3v1024x8m81_0/LWL[87] xdec128_3v1024x8m81_0/RWL[30] xdec128_3v1024x8m81_0/RWL[121]
+ xdec128_3v1024x8m81_0/LWL[83] xdec128_3v1024x8m81_0/LWL[51] xdec128_3v1024x8m81_0/LWL[46]
+ control_3v1024x8_3v1024x8m81_0/xc[3] xdec128_3v1024x8m81_0/LWL[104] xdec128_3v1024x8m81_0/RWL[26]
+ xdec128_3v1024x8m81_0/LWL[107] xdec128_3v1024x8m81_0/RWL[67] control_3v1024x8_3v1024x8m81_0/xc[2]
+ xdec128_3v1024x8m81_0/LWL[124] xdec128_3v1024x8m81_0/LWL[103] xdec128_3v1024x8m81_0/RWL[33]
+ xdec128_3v1024x8m81_0/LWL[11] xdec128_3v1024x8m81_0/LWL[70] xdec128_3v1024x8m81_0/LWL[18]
+ xdec128_3v1024x8m81_0/LWL[80] xdec128_3v1024x8m81_0/LWL[44] xdec128_3v1024x8m81_0/RWL[61]
+ xdec128_3v1024x8m81_0/RWL[104] xdec128_3v1024x8m81_0/LWL[90] xdec128_3v1024x8m81_0/RWL[24]
+ xdec128_3v1024x8m81_0/RWL[27] xdec128_3v1024x8m81_0/LWL[39] xdec128_3v1024x8m81_0/RWL[77]
+ xdec128_3v1024x8m81_0/RWL[114] xdec128_3v1024x8m81_0/RWL[34] xdec128_3v1024x8m81_0/LWL[4]
+ xdec128_3v1024x8m81_0/LWL[113] xdec128_3v1024x8m81_0/RWL[124] xdec128_3v1024x8m81_0/LWL[47]
+ xdec128_3v1024x8m81_0/RWL[16] xdec128_3v1024x8m81_0/LWL[23] xdec128_3v1024x8m81_0/RWL[70]
+ xdec128_3v1024x8m81_0/LWL[62] xdec128_3v1024x8m81_0/RWL[31] xdec128_3v1024x8m81_0/LWL[31]
+ xdec128_3v1024x8m81_0/RWL[41] xdec128_3v1024x8m81_0/RWL[80] xdec128_3v1024x8m81_0/LWL[42]
+ xdec128_3v1024x8m81_0/LWL[106] xdec128_3v1024x8m81_0/RWL[7] xdec128_3v1024x8m81_0/RWL[52]
+ xdec128_3v1024x8m81_0/RWL[22] xdec128_3v1024x8m81_0/LWL[7] xdec128_3v1024x8m81_0/LWL[127]
+ xdec128_3v1024x8m81_0/RWL[49] xdec128_3v1024x8m81_0/RWL[87] xdec128_3v1024x8m81_0/LWL[116]
+ VDD xdec128_3v1024x8m81_0/RWL[15] xdec128_3v1024x8m81_0/LWL[32] xdec128_3v1024x8m81_0/LWL[2]
+ xdec128_3v1024x8m81_0/LWL[126] xdec128_3v1024x8m81_0/LWL[123] xdec128_3v1024x8m81_0/RWL[14]
+ xdec128_3v1024x8m81_0/RWL[83] xdec128_3v1024x8m81_0/LWL[49] xdec128_3v1024x8m81_0/LWL[72]
+ xdec128_3v1024x8m81_0/LWL[60] xdec128_3v1024x8m81_0/RWL[107] VSS xdec128_3v1024x8m81
.ends

