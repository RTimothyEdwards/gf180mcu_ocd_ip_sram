magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< polysilicon >>
rect -14 1058 41 1092
rect -14 -34 41 0
use nmos_5p0431059130205_3v512x8m81  nmos_5p0431059130205_3v512x8m81_0
timestamp 1763765945
transform 1 0 -14 0 1 0
box -88 -44 144 1102
<< end >>
