magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< psubdiff >>
rect -1382 23 1382 56
rect -1382 -23 -1240 23
rect 1351 -23 1382 23
rect -1382 -56 1382 -23
<< psubdiffcont >>
rect -1240 -23 1351 23
<< metal1 >>
rect -1368 23 1368 41
rect -1368 -23 -1240 23
rect 1351 -23 1368 23
rect -1368 -42 1368 -23
<< end >>
