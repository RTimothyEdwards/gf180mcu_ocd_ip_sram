magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_0
array 0 7 -436 0 31 1212
timestamp 1763765945
transform -1 0 12924 0 1 0
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1
array 0 7 -436 0 31 1212
timestamp 1763765945
transform -1 0 5108 0 1 0
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_2
array 0 7 436 0 31 1212
timestamp 1763765945
transform 1 0 600 0 1 0
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_3
array 0 7 436 0 31 1212
timestamp 1763765945
transform 1 0 8416 0 1 0
box 62 103 538 1445
use 018SRAM_strap1_2x_512x8m81  018SRAM_strap1_2x_512x8m81_0
array 0 0 -420 0 31 1212
timestamp 1763765945
transform -1 0 12497 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_2x_512x8m81  018SRAM_strap1_2x_512x8m81_1
array 0 0 -420 0 31 1212
timestamp 1763765945
transform -1 0 773 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_2x_512x8m81  018SRAM_strap1_2x_512x8m81_2
array 0 0 -420 0 31 1212
timestamp 1763765945
transform -1 0 4681 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_2x_512x8m81  018SRAM_strap1_2x_512x8m81_3
array 0 0 -420 0 31 1212
timestamp 1763765945
transform -1 0 8589 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_2x_bndry_512x8m81  018SRAM_strap1_2x_bndry_512x8m81_0
array 0 0 420 0 31 1212
timestamp 1763765945
transform 1 0 15803 0 1 900
box 91 -797 511 545
<< end >>
