magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< error_p >>
rect -79 -8 -33 64
rect 126 -8 172 64
<< nmos >>
rect 0 0 93 56
<< ndiff >>
rect -92 56 -20 64
rect 113 56 185 64
rect -92 51 0 56
rect -92 5 -79 51
rect -33 5 0 51
rect -92 0 0 5
rect 93 51 185 56
rect 93 5 126 51
rect 172 5 185 51
rect 93 0 185 5
rect -92 -8 -20 0
rect 113 -8 185 0
<< ndiffc >>
rect -79 5 -33 51
rect 126 5 172 51
<< polysilicon >>
rect 0 56 93 100
rect 0 -44 93 0
<< metal1 >>
rect -79 51 -33 64
rect -79 -8 -33 5
rect 126 51 172 64
rect 126 -8 172 5
<< labels >>
flabel ndiffc -44 28 -44 28 0 FreeSans 93 0 0 0 S
flabel ndiffc 137 28 137 28 0 FreeSans 93 0 0 0 D
<< end >>
