magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect -133 -65 160 1589
<< polysilicon >>
rect -14 1523 41 1557
rect -14 -34 41 0
use pmos_5p04310591302070_512x8m81  pmos_5p04310591302070_512x8m81_0
timestamp 1763476864
transform 1 0 -14 0 1 0
box -174 -86 230 1610
<< end >>
