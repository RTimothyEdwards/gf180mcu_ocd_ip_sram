magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal2 >>
rect -119 172 119 198
rect -119 -132 -93 172
rect 93 -132 119 172
rect -119 -158 119 -132
<< via2 >>
rect -93 -132 93 172
<< metal3 >>
rect -119 172 119 198
rect -119 -132 -93 172
rect 93 -132 119 172
rect -119 -158 119 -132
<< end >>
