magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal1 >>
rect -44 26 635 46
rect -44 -26 -26 26
rect 617 -26 635 26
rect -44 -46 635 -26
<< via1 >>
rect -26 -26 617 26
<< metal2 >>
rect -45 26 635 46
rect -45 -26 -26 26
rect 617 -26 635 26
rect -45 -46 635 -26
<< end >>
