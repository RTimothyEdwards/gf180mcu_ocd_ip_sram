magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< error_s >>
rect -117 0 -71 106
rect 43 0 89 106
rect 203 0 249 106
<< polysilicon >>
rect -42 106 13 140
rect 118 106 174 140
rect -42 -34 13 0
rect 118 -34 174 0
use pmos_5p0431059130203_256x8m81  pmos_5p0431059130203_256x8m81_0
timestamp 1763766357
transform 1 0 -14 0 1 0
box -202 -86 362 192
<< end >>
