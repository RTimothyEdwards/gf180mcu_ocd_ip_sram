magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nmos >>
rect 0 0 56 149
<< ndiff >>
rect -88 135 0 149
rect -88 13 -75 135
rect -29 13 0 135
rect -88 0 0 13
rect 56 135 144 149
rect 56 13 85 135
rect 131 13 144 135
rect 56 0 144 13
<< ndiffc >>
rect -75 13 -29 135
rect 85 13 131 135
<< polysilicon >>
rect 0 149 56 193
rect 0 -44 56 0
<< metal1 >>
rect -75 135 -29 149
rect -75 0 -29 13
rect 85 135 131 149
rect 85 0 131 13
<< labels >>
flabel ndiffc -40 74 -40 74 0 FreeSans 93 0 0 0 S
flabel ndiffc 96 74 96 74 0 FreeSans 93 0 0 0 D
<< end >>
