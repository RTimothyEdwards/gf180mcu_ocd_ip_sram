magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal2 >>
rect -70 236 70 243
rect -70 -236 -63 236
rect 63 -236 70 236
rect -70 -243 70 -236
<< via2 >>
rect -63 -236 63 236
<< metal3 >>
rect -70 236 70 243
rect -70 -236 -63 236
rect 63 -236 70 236
rect -70 -243 70 -236
<< end >>
