magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal1 >>
rect -118 100 119 128
rect -118 -106 -92 100
rect -119 -170 -92 -106
rect 92 -170 119 100
rect -119 -198 119 -170
<< via1 >>
rect -92 -170 92 100
<< metal2 >>
rect -118 100 119 128
rect -118 -170 -92 100
rect 92 -170 119 100
rect -118 -198 119 -170
<< end >>
