magic
tech gf180mcuD
magscale 1 10
timestamp 1765833244
<< polysilicon >>
rect -289 23 289 48
rect -289 -23 -244 23
rect 244 -23 289 23
rect -289 -48 289 -23
<< polycontact >>
rect -244 -23 244 23
<< metal1 >>
rect -261 23 261 42
rect -261 -23 -244 23
rect 244 -23 261 23
rect -261 -42 261 -23
<< end >>
