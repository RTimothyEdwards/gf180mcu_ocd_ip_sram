* NGSPICE file created from gf180mcu_ocd_ip_sram__sram256x8m8wm1.ext - technology: gf180mcuD

.subckt x018SRAM_cell1_dummy_3v256x8m81 m3_82_330# a_248_342# a_248_592# w_82_512#
+ a_62_178# m2_346_89# m2_134_89# VSUBS
X0 a_248_592# a_192_298# a_110_250# w_82_512# pfet_03v3 ad=0.1613p pd=1.39u as=0.1238p ps=1.44u w=0.28u l=0.28u
X1 a_248_342# a_192_298# a_110_250# VSUBS nfet_03v3 ad=0.171p pd=1.33u as=0.15665p ps=1.32u w=0.45u l=0.28u
X2 a_192_298# a_110_250# a_248_592# w_82_512# pfet_03v3 ad=0.1238p pd=1.44u as=0.1613p ps=1.39u w=0.28u l=0.28u
X3 a_192_298# a_110_250# a_248_342# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.171p ps=1.33u w=0.45u l=0.28u
X4 a_110_250# a_62_178# a_110_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
X5 a_192_298# a_62_178# a_430_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
.ends

.subckt new_dummyrow_unit_3v256x8m81 018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89# 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89# VSUBS 018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89#
X018SRAM_cell1_dummy_3v256x8m81_10 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_11 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_12 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_13 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_15 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_14 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_0 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_1 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_2 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_3 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_4 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_5 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_6 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_7 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_8 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_9 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
.ends

.subckt new_dummyrowunit01_3v256x8m81 018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89#
+ VSUBS 018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89#
X018SRAM_cell1_dummy_3v256x8m81_10 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_11 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_12 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_13 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_15 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_14 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_0 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_1 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_2 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_3 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_4 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_5 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_6 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_7 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_8 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_9 018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS 018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
.ends

.subckt x018SRAM_cell1_3v256x8m81 m3_82_330# a_248_342# a_248_592# a_62_178# w_30_512#
+ a_430_96# a_110_96# VSUBS
X0 a_248_592# a_192_298# a_110_250# w_30_512# pfet_03v3 ad=0.1613p pd=1.39u as=0.1238p ps=1.44u w=0.28u l=0.28u
X1 a_248_342# a_192_298# a_110_250# VSUBS nfet_03v3 ad=0.171p pd=1.33u as=0.15665p ps=1.32u w=0.45u l=0.28u
X2 a_192_298# a_110_250# a_248_592# w_30_512# pfet_03v3 ad=0.1238p pd=1.44u as=0.1613p ps=1.39u w=0.28u l=0.28u
X3 a_192_298# a_110_250# a_248_342# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.171p ps=1.33u w=0.45u l=0.28u
X4 a_110_250# a_62_178# a_110_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
X5 a_192_298# a_62_178# a_430_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
.ends

.subckt x018SRAM_cell1_cutPC_3v256x8m81 m3_82_330# a_248_342# a_248_592# a_62_178#
+ w_30_512# a_430_96# a_110_96# VSUBS
X0 a_248_592# a_192_298# a_110_250# w_30_512# pfet_03v3 ad=0.1613p pd=1.39u as=0.1238p ps=1.44u w=0.28u l=0.28u
X1 a_248_342# a_192_298# a_110_250# VSUBS nfet_03v3 ad=0.171p pd=1.33u as=0.15665p ps=1.32u w=0.45u l=0.28u
X2 a_192_298# a_110_250# a_248_592# w_30_512# pfet_03v3 ad=0.1238p pd=1.44u as=0.1613p ps=1.39u w=0.28u l=0.28u
X3 a_192_298# a_110_250# a_248_342# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.171p ps=1.33u w=0.45u l=0.28u
X4 a_110_250# a_62_178# a_110_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
X5 a_192_298# a_62_178# a_430_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
.ends

.subckt array16_256_dummy_01_3v256x8m81 018SRAM_cell1_cutPC_3v256x8m81_55/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_10/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_10/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_51/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_51/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_2/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_53/a_248_592#
+ 018SRAM_cell1_cutPC_3v256x8m81_6/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_2/a_248_592#
+ 018SRAM_cell1_cutPC_3v256x8m81_50/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_11/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_11/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_2/w_30_512#
+ 018SRAM_cell1_cutPC_3v256x8m81_50/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_61/a_62_178#
+ VDD_uq0 018SRAM_cell1_cutPC_3v256x8m81_60/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_60/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_3/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_3/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_31/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_13/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_52/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_31/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_3/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_61/a_248_592#
+ 018SRAM_cell1_cutPC_3v256x8m81_51/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_51/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_12/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_12/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_7/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_61/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_61/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_4/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_4/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_51/a_248_592#
+ 018SRAM_cell1_cutPC_3v256x8m81_3/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_56/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_50/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_52/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_4/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_52/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_13/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_52/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_13/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_62/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_62/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_7/w_30_512#
+ 018SRAM_cell1_cutPC_3v256x8m81_5/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_5/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_50/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_3/w_30_512#
+ VSS_uq0 018SRAM_cell1_cutPC_3v256x8m81_5/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_62/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_53/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_14/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_53/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_14/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_14/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_63/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_63/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_6/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_6/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_10/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_49/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_8/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_6/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_54/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_15/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_15/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_54/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_4/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_62/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_57/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# 018SRAM_cell1_cutPC_3v256x8m81_7/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_0/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_7/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_49/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_48/a_248_592#
+ 018SRAM_cell1_cutPC_3v256x8m81_53/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_53/w_30_512#
+ 018SRAM_cell1_cutPC_3v256x8m81_7/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_55/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_55/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_8/w_30_512#
+ 018SRAM_cell1_cutPC_3v256x8m81_4/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_8/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_8/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_63/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_0/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_8/a_248_592#
+ 018SRAM_cell1_cutPC_3v256x8m81_48/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_15/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_56/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_56/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_11/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_9/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_9/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_5/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_58/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_57/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v256x8m81_57/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_54/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_48/w_30_512#
+ 018SRAM_cell1_cutPC_3v256x8m81_52/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_50/a_62_178#
+ VDD VSS 018SRAM_cell1_cutPC_3v256x8m81_48/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_48/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_58/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_5/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_58/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_31/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_0/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_60/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_49/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_49/m3_82_330#
+ 018SRAM_cell1_cutPC_3v256x8m81_49/a_248_342# 018SRAM_cell1_cutPC_3v256x8m81_12/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_59/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_59/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_61/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_6/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_59/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_2/a_62_178#
+ VSUBS
X018SRAM_cell1_cutPC_3v256x8m81_4 018SRAM_cell1_cutPC_3v256x8m81_4/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_4/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_4/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_4/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_4/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_5 018SRAM_cell1_cutPC_3v256x8m81_5/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_5/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_5/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_5/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_5/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_6 018SRAM_cell1_cutPC_3v256x8m81_6/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_6/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_6/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_6/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_6/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_8 018SRAM_cell1_cutPC_3v256x8m81_8/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_8/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_8/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_8/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_8/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_7 018SRAM_cell1_cutPC_3v256x8m81_7/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_7/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_7/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_7/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_7/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_9 018SRAM_cell1_cutPC_3v256x8m81_9/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_9/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_9/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_60 018SRAM_cell1_cutPC_3v256x8m81_60/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_60/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_3/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_60/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_3/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_50 018SRAM_cell1_cutPC_3v256x8m81_50/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_50/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_50/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_50/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_50/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_61 018SRAM_cell1_cutPC_3v256x8m81_61/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_61/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_61/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_61/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_61/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_51 018SRAM_cell1_cutPC_3v256x8m81_51/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_51/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_51/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_51/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_51/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_62 018SRAM_cell1_cutPC_3v256x8m81_62/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_62/a_248_342#
+ VDD_uq0 018SRAM_cell1_cutPC_3v256x8m81_62/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_62/w_30_512#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_52 018SRAM_cell1_cutPC_3v256x8m81_52/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_52/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_52/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_52/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_52/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_53 018SRAM_cell1_cutPC_3v256x8m81_53/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_53/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_53/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_53/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_53/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_31 018SRAM_cell1_cutPC_3v256x8m81_31/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_31/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_61/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_31/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_61/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_63 018SRAM_cell1_cutPC_3v256x8m81_63/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_63/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_2/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_63/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_2/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_10 018SRAM_cell1_cutPC_3v256x8m81_10/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_10/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_53/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_10/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_53/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_54 018SRAM_cell1_cutPC_3v256x8m81_54/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_54/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_54/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_11 018SRAM_cell1_cutPC_3v256x8m81_11/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_11/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_52/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_11/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_52/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_55 018SRAM_cell1_cutPC_3v256x8m81_55/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_55/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_8/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_55/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_8/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_12 018SRAM_cell1_cutPC_3v256x8m81_12/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_12/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_51/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_12/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_51/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_56 018SRAM_cell1_cutPC_3v256x8m81_56/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_56/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_7/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_56/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_7/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_13 018SRAM_cell1_cutPC_3v256x8m81_13/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_13/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_50/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_13/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_50/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_57 018SRAM_cell1_cutPC_3v256x8m81_57/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_57/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_6/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_57/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_6/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_14 018SRAM_cell1_cutPC_3v256x8m81_14/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_14/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_49/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_14/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_49/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_58 018SRAM_cell1_cutPC_3v256x8m81_58/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_58/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_5/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_58/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_5/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_48 018SRAM_cell1_cutPC_3v256x8m81_48/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_48/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_48/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_48/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_48/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_15 018SRAM_cell1_cutPC_3v256x8m81_15/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_15/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_48/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_15/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_48/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_59 018SRAM_cell1_cutPC_3v256x8m81_59/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_59/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_4/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_59/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_4/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_49 018SRAM_cell1_cutPC_3v256x8m81_49/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_49/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_49/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_49/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_49/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_0 018SRAM_cell1_cutPC_3v256x8m81_0/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_0/a_248_342#
+ VDD 018SRAM_cell1_cutPC_3v256x8m81_0/a_62_178# 018SRAM_cell1_cutPC_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96# 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96#
+ VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_2 018SRAM_cell1_cutPC_3v256x8m81_2/m3_82_330# VSS_uq0
+ 018SRAM_cell1_cutPC_3v256x8m81_2/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_2/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_2/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
X018SRAM_cell1_cutPC_3v256x8m81_3 018SRAM_cell1_cutPC_3v256x8m81_3/m3_82_330# 018SRAM_cell1_cutPC_3v256x8m81_3/a_248_342#
+ 018SRAM_cell1_cutPC_3v256x8m81_3/a_248_592# 018SRAM_cell1_cutPC_3v256x8m81_3/a_62_178#
+ 018SRAM_cell1_cutPC_3v256x8m81_3/w_30_512# 018SRAM_cell1_cutPC_3v256x8m81_9/a_430_96#
+ 018SRAM_cell1_cutPC_3v256x8m81_9/a_110_96# VSUBS x018SRAM_cell1_cutPC_3v256x8m81
.ends

.subckt ldummy_3v256x4_3v256x8m81 array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_3/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_53/a_248_592# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_3/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_23/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_23/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_3/a_248_592#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_11/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_7/w_30_512#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_50/m3_82_330# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_11/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_50/a_248_342# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_3/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_60/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_60/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_4/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_31/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_52/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_31/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_4/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_24/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_24/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_50/w_30_512# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_4/a_248_592# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_51/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_61/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_12/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_12/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_51/a_248_342# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_61/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_61/a_248_342#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_5/m3_82_330# 018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_5/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_51/a_248_592#
+ 018SRAM_cell1_dummy_3v256x8m81_25/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_25/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_5/a_248_592#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_52/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_13/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_52/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_13/a_248_342# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_62/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/VSS_uq0 array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_62/a_248_342#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_16/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_16/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_6/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_6/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_50/a_248_592# 018SRAM_cell1_dummy_3v256x8m81_26/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_26/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_8/w_30_512#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_6/a_248_592# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_4/w_30_512#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_53/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_14/m3_82_330#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_53/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_14/a_248_342# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_63/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_63/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_17/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_17/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_7/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_7/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_49/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_49/a_248_592#
+ 018SRAM_cell1_dummy_3v256x8m81_27/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_27/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_53/w_30_512#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_7/a_248_592# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_54/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_15/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_15/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_54/a_248_342#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_18/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_18/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_8/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_8/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_48/a_248_592# 018SRAM_cell1_dummy_3v256x8m81_28/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_28/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_8/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_55/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_55/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_19/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_9/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_19/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_9/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_9/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_5/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_29/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_29/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_9/a_248_592# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_56/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_56/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_48/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_52/w_30_512# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_57/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_57/m3_82_330# 018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_0/m3_82_330# 018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_0/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_20/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_20/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_48/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_30/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_48/a_248_342# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_30/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_58/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_58/a_248_342# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_6/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_61/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_2/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_21/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_21/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_49/m3_82_330# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_49/a_248_342# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_31/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_31/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_59/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_59/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_51/w_30_512# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_2/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_22/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_22/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89# array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_2/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_10/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_10/a_248_342#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89#
+ VSUBS 018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ array16_256_dummy_01_3v256x8m81_0/VDD new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89#
Xnew_dummyrow_unit_3v256x8m81_0 new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ array16_256_dummy_01_3v256x8m81_0/VDD new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89#
+ VSUBS new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ VSUBS new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# new_dummyrow_unit_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89#
+ new_dummyrow_unit_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_10 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_21 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_21/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_21/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_11 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_22 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_22/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_22/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_12 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_23 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_23/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_23/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_13 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_24 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_24/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_24/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_14 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_25 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_25/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_25/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_26 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_26/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_26/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_15 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_16 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_16/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_16/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_27 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_27/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_27/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_17 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_17/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_17/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_28 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_28/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_28/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_18 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_18/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_18/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_29 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_29/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_29/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_19 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_19/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_19/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
Xnew_dummyrowunit01_3v256x8m81_0 new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89#
+ array16_256_dummy_01_3v256x8m81_0/VDD VSUBS new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89#
+ VSUBS new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ new_dummyrowunit01_3v256x8m81_0/018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89# new_dummyrowunit01_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_0 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_3v256x8m81_0 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0 018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# VSUBS x018SRAM_cell1_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_1 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_3v256x8m81_1 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD VSUBS
+ array16_256_dummy_01_3v256x8m81_0/VDD 018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_3v256x8m81_1/a_110_96#
+ VSUBS x018SRAM_cell1_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_2 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_3 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_4 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_5 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
Xarray16_256_dummy_01_3v256x8m81_0 VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_10/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_10/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_51/w_30_512#
+ VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_2/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_53/a_248_592# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_6/w_30_512#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_2/a_248_592# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_50/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_11/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_11/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_2/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_50/a_248_342#
+ VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0 array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_60/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_60/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_3/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_3/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_31/m3_82_330#
+ VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_52/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_31/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_3/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_61/a_248_592# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_51/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_51/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_12/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_12/m3_82_330# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_61/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_61/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_4/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_4/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_51/a_248_592# VSUBS
+ VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_50/w_30_512#
+ VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_4/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_52/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_13/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_52/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_13/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_62/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_62/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_7/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_5/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_5/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_50/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_3/w_30_512# array16_256_dummy_01_3v256x8m81_0/VSS_uq0
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_5/a_248_592# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_53/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_14/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_53/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_14/a_248_342#
+ VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_63/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_63/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_6/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_6/a_248_342# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_49/a_248_592# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_6/a_248_592# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_54/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_15/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_15/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_54/a_248_342# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_3v256x8m81_1/a_110_96#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_7/a_248_342# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_7/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_49/w_30_512#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_48/a_248_592# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_53/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_7/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_55/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_55/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_8/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_4/w_30_512#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_8/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_8/m3_82_330#
+ VSUBS array16_256_dummy_01_3v256x8m81_0/VDD array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_8/a_248_592#
+ VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_56/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_56/m3_82_330# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_9/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_9/a_248_342#
+ VSUBS VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_9/a_248_592#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_57/m3_82_330# 018SRAM_cell1_3v256x8m81_1/a_430_96#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_57/a_248_342# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_48/w_30_512# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_52/w_30_512#
+ VSUBS array16_256_dummy_01_3v256x8m81_0/VDD VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_48/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_48/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_9/w_30_512#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_58/a_248_342# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_5/w_30_512#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_58/m3_82_330# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_0/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_0/a_248_342#
+ VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_49/m3_82_330#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_49/a_248_342# VSUBS
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_59/m3_82_330# array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_59/a_248_342#
+ array16_256_dummy_01_3v256x8m81_0/018SRAM_cell1_cutPC_3v256x8m81_61/w_30_512# VSUBS
+ VSUBS VSUBS VSUBS array16_256_dummy_01_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_6 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_7 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_9 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_8 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_30 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_30/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_30/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_31 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_31/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_31/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_20 VSUBS VSUBS array16_256_dummy_01_3v256x8m81_0/VDD_uq0
+ array16_256_dummy_01_3v256x8m81_0/VDD_uq0 VSUBS 018SRAM_cell1_dummy_3v256x8m81_20/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_20/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
.ends

.subckt pmos_5p04310591302030_3v256x8m81 D_uq2 a_871_n45# D_uq1 D_uq0 D a_n252_n45#
+ a_550_n45# a_229_n45# w_n426_n86# S_uq4 S_uq2 S_uq3 S_uq1 S_uq0 a_390_n45# S a_n92_n45#
+ a_1032_n45# a_1192_n45# D_uq3 a_711_n45# a_69_n45#
X0 D_uq1 a_390_n45# S_uq2 w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.33205p ps=1.79u w=1.265u l=0.28u
X1 D_uq3 a_n252_n45# S_uq4 w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.5566p ps=3.41u w=1.265u l=0.28u
X2 D_uq2 a_69_n45# S_uq3 w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.33205p ps=1.79u w=1.265u l=0.28u
X3 S_uq2 a_229_n45# D_uq2 w_n426_n86# pfet_03v3 ad=0.33205p pd=1.79u as=0.3289p ps=1.785u w=1.265u l=0.28u
X4 S_uq1 a_550_n45# D_uq1 w_n426_n86# pfet_03v3 ad=0.33205p pd=1.79u as=0.3289p ps=1.785u w=1.265u l=0.28u
X5 S_uq0 a_1192_n45# D_uq0 w_n426_n86# pfet_03v3 ad=0.5566p pd=3.41u as=0.3289p ps=1.785u w=1.265u l=0.28u
X6 D_uq0 a_1032_n45# S w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.33205p ps=1.79u w=1.265u l=0.28u
X7 S_uq3 a_n92_n45# D_uq3 w_n426_n86# pfet_03v3 ad=0.33205p pd=1.79u as=0.3289p ps=1.785u w=1.265u l=0.28u
X8 S a_871_n45# D w_n426_n86# pfet_03v3 ad=0.33205p pd=1.79u as=0.3289p ps=1.785u w=1.265u l=0.28u
X9 D a_711_n45# S_uq1 w_n426_n86# pfet_03v3 ad=0.3289p pd=1.785u as=0.33205p ps=1.79u w=1.265u l=0.28u
.ends

.subckt pmos_1p2$$45095980_3v256x8m81 a_697_n34# pmos_5p04310591302030_3v256x8m81_0/D
+ a_n106_n34# a_n266_n34# pmos_5p04310591302030_3v256x8m81_0/S_uq4 a_376_n34# pmos_5p04310591302030_3v256x8m81_0/S_uq3
+ pmos_5p04310591302030_3v256x8m81_0/S_uq2 pmos_5p04310591302030_3v256x8m81_0/S_uq0
+ pmos_5p04310591302030_3v256x8m81_0/S_uq1 a_1018_n34# a_1178_n34# a_55_n34# a_857_n34#
+ pmos_5p04310591302030_3v256x8m81_0/D_uq2 pmos_5p04310591302030_3v256x8m81_0/D_uq3
+ pmos_5p04310591302030_3v256x8m81_0/D_uq1 pmos_5p04310591302030_3v256x8m81_0/D_uq0
+ pmos_5p04310591302030_3v256x8m81_0/S a_536_n34# w_987_n66# a_215_n34#
Xpmos_5p04310591302030_3v256x8m81_0 pmos_5p04310591302030_3v256x8m81_0/D_uq2 a_857_n34#
+ pmos_5p04310591302030_3v256x8m81_0/D_uq1 pmos_5p04310591302030_3v256x8m81_0/D_uq0
+ pmos_5p04310591302030_3v256x8m81_0/D a_n266_n34# a_536_n34# a_215_n34# w_987_n66#
+ pmos_5p04310591302030_3v256x8m81_0/S_uq4 pmos_5p04310591302030_3v256x8m81_0/S_uq2
+ pmos_5p04310591302030_3v256x8m81_0/S_uq3 pmos_5p04310591302030_3v256x8m81_0/S_uq1
+ pmos_5p04310591302030_3v256x8m81_0/S_uq0 a_376_n34# pmos_5p04310591302030_3v256x8m81_0/S
+ a_n106_n34# a_1018_n34# a_1178_n34# pmos_5p04310591302030_3v256x8m81_0/D_uq3 a_697_n34#
+ a_55_n34# pmos_5p04310591302030_3v256x8m81
.ends

.subckt pmos_5p04310591302027_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.28u
.ends

.subckt pmos_5p04310591302024_3v256x8m81 w_n286_n86# D_uq1 D_uq0 a_530_n44# D a_n112_n44#
+ a_209_n44# a_369_n44# a_48_n44# S_uq1 S_uq0 S
X0 D_uq1 a_n112_n44# S_uq1 w_n286_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X1 S_uq0 a_369_n44# D w_n286_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D a_209_n44# S w_n286_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.27692p ps=1.58u w=1.055u l=0.28u
X3 D_uq0 a_530_n44# S_uq0 w_n286_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.27692p ps=1.58u w=1.055u l=0.28u
X4 S a_48_n44# D_uq1 w_n286_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46282796_3v256x8m81 pmos_5p04310591302024_3v256x8m81_0/S a_n126_n34#
+ pmos_5p04310591302024_3v256x8m81_0/S_uq1 pmos_5p04310591302024_3v256x8m81_0/S_uq0
+ a_195_n34# pmos_5p04310591302024_3v256x8m81_0/D pmos_5p04310591302024_3v256x8m81_0/D_uq1
+ a_516_n34# pmos_5p04310591302024_3v256x8m81_0/D_uq0 w_163_n66# a_355_n34# a_34_n34#
Xpmos_5p04310591302024_3v256x8m81_0 w_163_n66# pmos_5p04310591302024_3v256x8m81_0/D_uq1
+ pmos_5p04310591302024_3v256x8m81_0/D_uq0 a_516_n34# pmos_5p04310591302024_3v256x8m81_0/D
+ a_n126_n34# a_195_n34# a_355_n34# a_34_n34# pmos_5p04310591302024_3v256x8m81_0/S_uq1
+ pmos_5p04310591302024_3v256x8m81_0/S_uq0 pmos_5p04310591302024_3v256x8m81_0/S pmos_5p04310591302024_3v256x8m81
.ends

.subckt nmos_5p04310591302029_3v256x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.54067p pd=3.32u as=0.3159p ps=1.735u w=1.215u l=0.28u
.ends

.subckt nmos_1p2$$45100076_3v256x8m81 nmos_5p04310591302029_3v256x8m81_0/S nmos_5p04310591302029_3v256x8m81_0/D
+ a_118_n34# a_n41_n34# nmos_5p04310591302029_3v256x8m81_0/S_uq0 VSUBS
Xnmos_5p04310591302029_3v256x8m81_0 nmos_5p04310591302029_3v256x8m81_0/D a_n41_n34#
+ a_118_n34# nmos_5p04310591302029_3v256x8m81_0/S_uq0 nmos_5p04310591302029_3v256x8m81_0/S
+ VSUBS nmos_5p04310591302029_3v256x8m81
.ends

.subckt nmos_5p04310591302032_3v256x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.1378p pd=1.05u as=0.2332p ps=1.94u w=0.53u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.23585p pd=1.95u as=0.1378p ps=1.05u w=0.53u l=0.28u
.ends

.subckt pmos_5p04310591302022_3v256x8m81 D_uq2 D_uq1 D_uq0 D a_n252_n44# a_550_n44#
+ a_229_n44# w_n426_n86# S_uq4 S_uq2 S_uq3 S_uq1 a_390_n44# S_uq0 S a_n92_n44# a_1032_n44#
+ a_1192_n44# a_711_n44# a_69_n44# D_uq3 a_871_n44#
X0 D_uq1 a_390_n44# S_uq2 w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.50005p ps=2.43u w=1.905u l=0.28u
X1 D_uq3 a_n252_n44# S_uq4 w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.8382p ps=4.69u w=1.905u l=0.28u
X2 D_uq2 a_69_n44# S_uq3 w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.50005p ps=2.43u w=1.905u l=0.28u
X3 S_uq2 a_229_n44# D_uq2 w_n426_n86# pfet_03v3 ad=0.50005p pd=2.43u as=0.4953p ps=2.425u w=1.905u l=0.28u
X4 S_uq1 a_550_n44# D_uq1 w_n426_n86# pfet_03v3 ad=0.50005p pd=2.43u as=0.4953p ps=2.425u w=1.905u l=0.28u
X5 S_uq0 a_1192_n44# D_uq0 w_n426_n86# pfet_03v3 ad=0.8382p pd=4.69u as=0.4953p ps=2.425u w=1.905u l=0.28u
X6 D_uq0 a_1032_n44# S w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.50005p ps=2.43u w=1.905u l=0.28u
X7 S_uq3 a_n92_n44# D_uq3 w_n426_n86# pfet_03v3 ad=0.50005p pd=2.43u as=0.4953p ps=2.425u w=1.905u l=0.28u
X8 S a_871_n44# D w_n426_n86# pfet_03v3 ad=0.50005p pd=2.43u as=0.4953p ps=2.425u w=1.905u l=0.28u
X9 D a_711_n44# S_uq1 w_n426_n86# pfet_03v3 ad=0.4953p pd=2.425u as=0.50005p ps=2.43u w=1.905u l=0.28u
.ends

.subckt pmos_1p2$$46283820_3v256x8m81 a_536_n34# pmos_5p04310591302022_3v256x8m81_0/D_uq3
+ pmos_5p04310591302022_3v256x8m81_0/D_uq2 a_215_n34# pmos_5p04310591302022_3v256x8m81_0/D_uq1
+ pmos_5p04310591302022_3v256x8m81_0/D_uq0 a_697_n34# a_n106_n34# a_n266_n34# pmos_5p04310591302022_3v256x8m81_0/S
+ a_376_n34# w_984_n66# a_1018_n34# a_1178_n34# pmos_5p04310591302022_3v256x8m81_0/S_uq4
+ pmos_5p04310591302022_3v256x8m81_0/S_uq3 a_55_n34# pmos_5p04310591302022_3v256x8m81_0/S_uq1
+ pmos_5p04310591302022_3v256x8m81_0/S_uq2 pmos_5p04310591302022_3v256x8m81_0/S_uq0
+ a_857_n34# pmos_5p04310591302022_3v256x8m81_0/D
Xpmos_5p04310591302022_3v256x8m81_0 pmos_5p04310591302022_3v256x8m81_0/D_uq2 pmos_5p04310591302022_3v256x8m81_0/D_uq1
+ pmos_5p04310591302022_3v256x8m81_0/D_uq0 pmos_5p04310591302022_3v256x8m81_0/D a_n266_n34#
+ a_536_n34# a_215_n34# w_984_n66# pmos_5p04310591302022_3v256x8m81_0/S_uq4 pmos_5p04310591302022_3v256x8m81_0/S_uq2
+ pmos_5p04310591302022_3v256x8m81_0/S_uq3 pmos_5p04310591302022_3v256x8m81_0/S_uq1
+ a_376_n34# pmos_5p04310591302022_3v256x8m81_0/S_uq0 pmos_5p04310591302022_3v256x8m81_0/S
+ a_n106_n34# a_1018_n34# a_1178_n34# a_697_n34# a_55_n34# pmos_5p04310591302022_3v256x8m81_0/D_uq3
+ a_857_n34# pmos_5p04310591302022_3v256x8m81
.ends

.subckt nmos_5p04310591302036_3v256x8m81 D_uq1 D_uq0 a_530_n44# D a_n112_n44# a_209_n44#
+ a_369_n44# a_48_n44# S_uq1 S_uq0 S VSUBS
X0 D_uq1 a_n112_n44# S_uq1 VSUBS nfet_03v3 ad=0.1378p pd=1.05u as=0.2332p ps=1.94u w=0.53u l=0.28u
X1 S_uq0 a_369_n44# D VSUBS nfet_03v3 ad=0.13913p pd=1.055u as=0.1378p ps=1.05u w=0.53u l=0.28u
X2 D a_209_n44# S VSUBS nfet_03v3 ad=0.1378p pd=1.05u as=0.13913p ps=1.055u w=0.53u l=0.28u
X3 D_uq0 a_530_n44# S_uq0 VSUBS nfet_03v3 ad=0.2332p pd=1.94u as=0.13913p ps=1.055u w=0.53u l=0.28u
X4 S a_48_n44# D_uq1 VSUBS nfet_03v3 ad=0.13913p pd=1.055u as=0.1378p ps=1.05u w=0.53u l=0.28u
.ends

.subckt nmos_1p2$$45101100_3v256x8m81 a_195_n34# nmos_5p04310591302036_3v256x8m81_0/S
+ a_35_n34# nmos_5p04310591302036_3v256x8m81_0/S_uq1 nmos_5p04310591302036_3v256x8m81_0/S_uq0
+ a_516_n34# nmos_5p04310591302036_3v256x8m81_0/D a_n125_n34# nmos_5p04310591302036_3v256x8m81_0/D_uq1
+ nmos_5p04310591302036_3v256x8m81_0/D_uq0 a_356_n34# VSUBS
Xnmos_5p04310591302036_3v256x8m81_0 nmos_5p04310591302036_3v256x8m81_0/D_uq1 nmos_5p04310591302036_3v256x8m81_0/D_uq0
+ a_516_n34# nmos_5p04310591302036_3v256x8m81_0/D a_n125_n34# a_195_n34# a_356_n34#
+ a_35_n34# nmos_5p04310591302036_3v256x8m81_0/S_uq1 nmos_5p04310591302036_3v256x8m81_0/S_uq0
+ nmos_5p04310591302036_3v256x8m81_0/S VSUBS nmos_5p04310591302036_3v256x8m81
.ends

.subckt nmos_5p04310591302033_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1576p pd=1.64u as=0.1576p ps=1.64u w=0.28u l=0.28u
.ends

.subckt pmos_5p04310591302031_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.4134p pd=2.11u as=0.6996p ps=4.06u w=1.59u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.6996p pd=4.06u as=0.4134p ps=2.11u w=1.59u l=0.28u
.ends

.subckt pmos_1p2$$46287916_3v256x8m81 w_n133_n66# pmos_5p04310591302031_3v256x8m81_0/S
+ a_n42_n34# pmos_5p04310591302031_3v256x8m81_0/D pmos_5p04310591302031_3v256x8m81_0/S_uq0
+ a_118_n34#
Xpmos_5p04310591302031_3v256x8m81_0 pmos_5p04310591302031_3v256x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302031_3v256x8m81_0/S_uq0 pmos_5p04310591302031_3v256x8m81_0/S
+ pmos_5p04310591302031_3v256x8m81
.ends

.subckt nmos_5p04310591302034_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.2948p pd=2.22u as=0.2948p ps=2.22u w=0.67u l=0.28u
.ends

.subckt pmos_5p04310591302035_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.2067p pd=1.315u as=0.3498p ps=2.47u w=0.795u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.3498p pd=2.47u as=0.2067p ps=1.315u w=0.795u l=0.28u
.ends

.subckt pmos_1p2$$46284844_3v256x8m81 w_n133_n66# pmos_5p04310591302035_3v256x8m81_0/S
+ pmos_5p04310591302035_3v256x8m81_0/S_uq0 pmos_5p04310591302035_3v256x8m81_0/D a_118_n34#
+ a_n42_n34#
Xpmos_5p04310591302035_3v256x8m81_0 pmos_5p04310591302035_3v256x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302035_3v256x8m81_0/S_uq0 pmos_5p04310591302035_3v256x8m81_0/S
+ pmos_5p04310591302035_3v256x8m81
.ends

.subckt nmos_5p04310591302026_3v256x8m81 D_uq2 D_uq1 D_uq0 a_154_n44# D a_n168_n44#
+ a_476_n44# a_798_n44# a_314_n44# S_uq2 S_uq1 a_n8_n44# S_uq0 S a_636_n44# VSUBS
X0 S_uq0 a_636_n44# D VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
X1 S a_314_n44# D_uq1 VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D_uq2 a_n168_n44# S_uq2 VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X3 S_uq1 a_n8_n44# D_uq2 VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
X4 D_uq0 a_798_n44# S_uq0 VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.27957p ps=1.585u w=1.055u l=0.28u
X5 D a_476_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.27957p ps=1.585u w=1.055u l=0.28u
X6 D_uq1 a_154_n44# S_uq1 VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.27957p ps=1.585u w=1.055u l=0.28u
.ends

.subckt nmos_1p2$$45102124_3v256x8m81 a_140_n34# nmos_5p04310591302026_3v256x8m81_0/S
+ a_462_n34# nmos_5p04310591302026_3v256x8m81_0/S_uq2 nmos_5p04310591302026_3v256x8m81_0/S_uq1
+ nmos_5p04310591302026_3v256x8m81_0/S_uq0 a_n181_n34# a_784_n34# a_300_n34# nmos_5p04310591302026_3v256x8m81_0/D
+ nmos_5p04310591302026_3v256x8m81_0/D_uq2 nmos_5p04310591302026_3v256x8m81_0/D_uq1
+ a_622_n34# a_n22_n34# nmos_5p04310591302026_3v256x8m81_0/D_uq0 VSUBS
Xnmos_5p04310591302026_3v256x8m81_0 nmos_5p04310591302026_3v256x8m81_0/D_uq2 nmos_5p04310591302026_3v256x8m81_0/D_uq1
+ nmos_5p04310591302026_3v256x8m81_0/D_uq0 a_140_n34# nmos_5p04310591302026_3v256x8m81_0/D
+ a_n181_n34# a_462_n34# a_784_n34# a_300_n34# nmos_5p04310591302026_3v256x8m81_0/S_uq2
+ nmos_5p04310591302026_3v256x8m81_0/S_uq1 a_n22_n34# nmos_5p04310591302026_3v256x8m81_0/S_uq0
+ nmos_5p04310591302026_3v256x8m81_0/S a_622_n34# VSUBS nmos_5p04310591302026_3v256x8m81
.ends

.subckt pmos_5p04310591302013_3v256x8m81 D_uq0 D a_265_n44# S_uq0 S a_n56_n44# a_104_n44#
+ w_n230_n86#
X0 D_uq0 a_265_n44# S_uq0 w_n230_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.27692p ps=1.58u w=1.055u l=0.28u
X1 D a_n56_n44# S w_n230_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X2 S_uq0 a_104_n44# D w_n230_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46286892_3v256x8m81 w_n133_n66# pmos_5p04310591302013_3v256x8m81_0/S_uq0
+ pmos_5p04310591302013_3v256x8m81_0/D pmos_5p04310591302013_3v256x8m81_0/D_uq0 a_251_n34#
+ a_n70_n34# a_90_n34# pmos_5p04310591302013_3v256x8m81_0/S
Xpmos_5p04310591302013_3v256x8m81_0 pmos_5p04310591302013_3v256x8m81_0/D_uq0 pmos_5p04310591302013_3v256x8m81_0/D
+ a_251_n34# pmos_5p04310591302013_3v256x8m81_0/S_uq0 pmos_5p04310591302013_3v256x8m81_0/S
+ a_n70_n34# a_90_n34# w_n133_n66# pmos_5p04310591302013_3v256x8m81
.ends

.subckt nmos_5p04310591302023_3v256x8m81 D a_n32_n44# a_136_n44# S_uq0 S VSUBS
X0 D a_n32_n44# S VSUBS nfet_03v3 ad=92.8f pd=0.92u as=0.1576p ps=1.64u w=0.28u l=0.28u
X1 S_uq0 a_136_n44# D VSUBS nfet_03v3 ad=0.159p pd=1.65u as=92.8f ps=0.92u w=0.28u l=0.28u
.ends

.subckt nmos_5p04310591302028_3v256x8m81 D_uq1 D_uq0 D a_64_n44# a_226_n44# a_386_n44#
+ a_548_n44# S_uq1 S_uq0 S a_n96_n44# VSUBS
X0 D_uq0 a_548_n44# S_uq0 VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.27957p ps=1.585u w=1.055u l=0.28u
X1 S_uq0 a_386_n44# D VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D a_226_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.27957p ps=1.585u w=1.055u l=0.28u
X3 D_uq1 a_n96_n44# S_uq1 VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X4 S a_64_n44# D_uq1 VSUBS nfet_03v3 ad=0.27957p pd=1.585u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_5p04310591302025_3v256x8m81 D_uq0 D a_265_n44# S_uq0 S a_n56_n44# a_104_n44#
+ w_n230_n85#
X0 D_uq0 a_265_n44# S_uq0 w_n230_n85# pfet_03v3 ad=0.9306p pd=5.11u as=0.55518p ps=2.64u w=2.115u l=0.28u
X1 D a_n56_n44# S w_n230_n85# pfet_03v3 ad=0.5499p pd=2.635u as=0.9306p ps=5.11u w=2.115u l=0.28u
X2 S_uq0 a_104_n44# D w_n230_n85# pfet_03v3 ad=0.55518p pd=2.64u as=0.5499p ps=2.635u w=2.115u l=0.28u
.ends

.subckt pmos_1p2$$46281772_3v256x8m81 pmos_5p04310591302025_3v256x8m81_0/S_uq0 pmos_5p04310591302025_3v256x8m81_0/S
+ a_251_n34# w_n133_n66# a_n70_n34# pmos_5p04310591302025_3v256x8m81_0/D_uq0 pmos_5p04310591302025_3v256x8m81_0/D
+ a_90_n34#
Xpmos_5p04310591302025_3v256x8m81_0 pmos_5p04310591302025_3v256x8m81_0/D_uq0 pmos_5p04310591302025_3v256x8m81_0/D
+ a_251_n34# pmos_5p04310591302025_3v256x8m81_0/S_uq0 pmos_5p04310591302025_3v256x8m81_0/S
+ a_n70_n34# a_90_n34# w_n133_n66# pmos_5p04310591302025_3v256x8m81
.ends

.subckt pmos_5p04310591302014_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.4642p ps=2.99u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46285868_3v256x8m81 w_n133_n66# pmos_5p04310591302014_3v256x8m81_0/S
+ pmos_5p04310591302014_3v256x8m81_0/D a_n14_n34#
Xpmos_5p04310591302014_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302014_3v256x8m81_0/S pmos_5p04310591302014_3v256x8m81
.ends

.subckt pmos_5p04310591302038_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.2464p pd=2u as=0.2464p ps=2u w=0.56u l=0.28u
.ends

.subckt nmos_5p04310591302037_3v256x8m81 a_20_n44# D a_181_n44# a_502_n44# S_uq2 a_662_n44#
+ a_n140_n44# S_uq0 a_341_n44# VSUBS
X0 S a_341_n44# D VSUBS nfet_03v3 ad=0.34912p pd=1.855u as=0.3458p ps=1.85u w=1.33u l=0.28u
X1 S_uq0 a_662_n44# D_uq0 VSUBS nfet_03v3 ad=0.5852p pd=3.54u as=0.3458p ps=1.85u w=1.33u l=0.28u
X2 D_uq0 a_502_n44# S VSUBS nfet_03v3 ad=0.3458p pd=1.85u as=0.34912p ps=1.855u w=1.33u l=0.28u
X3 S_uq1 a_20_n44# D_uq1 VSUBS nfet_03v3 ad=0.34912p pd=1.855u as=0.3458p ps=1.85u w=1.33u l=0.28u
X4 D a_181_n44# S_uq1 VSUBS nfet_03v3 ad=0.3458p pd=1.85u as=0.34912p ps=1.855u w=1.33u l=0.28u
X5 D_uq1 a_n140_n44# S_uq2 VSUBS nfet_03v3 ad=0.3458p pd=1.85u as=0.5852p ps=3.54u w=1.33u l=0.28u
.ends

.subckt nmos_1p2$$45103148_3v256x8m81 a_327_n34# a_n153_n34# a_488_n34# nmos_5p04310591302037_3v256x8m81_0/S_uq2
+ nmos_5p04310591302037_3v256x8m81_0/S_uq0 a_167_n34# a_6_n34# nmos_5p04310591302037_3v256x8m81_0/D
+ a_648_n34# VSUBS
Xnmos_5p04310591302037_3v256x8m81_0 a_6_n34# nmos_5p04310591302037_3v256x8m81_0/D
+ a_167_n34# a_488_n34# nmos_5p04310591302037_3v256x8m81_0/S_uq2 a_648_n34# a_n153_n34#
+ nmos_5p04310591302037_3v256x8m81_0/S_uq0 a_327_n34# VSUBS nmos_5p04310591302037_3v256x8m81
.ends

.subckt nmos_5p04310591302012_3v256x8m81 a_n83_n44# D_uq0 D a_77_n44# S_uq1 S_uq0
+ S a_237_n44# a_397_n44# VSUBS
X0 S a_77_n44# D VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.2743p ps=1.575u w=1.055u l=0.28u
X1 S_uq0 a_397_n44# D_uq0 VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D_uq0 a_237_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.2743p ps=1.575u w=1.055u l=0.28u
X3 D a_n83_n44# S_uq1 VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
.ends

.subckt sacntl_2_3v256x8m81 pcb se vdd_uq0 pmos_5p04310591302027_3v256x8m81_1/S_uq0
+ pmos_5p04310591302027_3v256x8m81_2/S_uq0 men vdd vss
Xpmos_1p2$$45095980_3v256x8m81_0 nmos_5p04310591302028_3v256x8m81_1/S se nmos_5p04310591302028_3v256x8m81_1/S
+ nmos_5p04310591302028_3v256x8m81_1/S vdd nmos_5p04310591302028_3v256x8m81_1/S vdd
+ vdd vdd vdd nmos_5p04310591302028_3v256x8m81_1/S nmos_5p04310591302028_3v256x8m81_1/S
+ nmos_5p04310591302028_3v256x8m81_1/S nmos_5p04310591302028_3v256x8m81_1/S se se
+ se se vdd nmos_5p04310591302028_3v256x8m81_1/S vdd nmos_5p04310591302028_3v256x8m81_1/S
+ pmos_1p2$$45095980_3v256x8m81
Xpmos_5p04310591302027_3v256x8m81_0 vdd_uq0 pmos_5p04310591302027_3v256x8m81_2/S_uq0
+ pmos_5p04310591302027_3v256x8m81_0/S vdd_uq0 pmos_5p04310591302027_3v256x8m81_0/S_uq0
+ pmos_5p04310591302027_3v256x8m81_0/S pmos_5p04310591302027_3v256x8m81
Xpmos_1p2$$46282796_3v256x8m81_0 vdd_uq0 men vdd_uq0 vdd_uq0 men pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D men pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ vdd_uq0 men men pmos_1p2$$46282796_3v256x8m81
Xpmos_5p04310591302027_3v256x8m81_1 vdd_uq0 pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ vss vdd_uq0 pmos_5p04310591302027_3v256x8m81_1/S_uq0 pmos_5p04310591302027_3v256x8m81_1/S
+ pmos_5p04310591302027_3v256x8m81
Xnmos_1p2$$45100076_3v256x8m81_0 vss pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ pmos_1p2$$46281772_3v256x8m81_1/pmos_5p04310591302025_3v256x8m81_0/S pmos_1p2$$46281772_3v256x8m81_1/pmos_5p04310591302025_3v256x8m81_0/S
+ vss vss nmos_1p2$$45100076_3v256x8m81
Xpmos_5p04310591302027_3v256x8m81_2 vdd_uq0 pmos_5p04310591302027_3v256x8m81_1/S_uq0
+ pmos_5p04310591302027_3v256x8m81_2/S vdd_uq0 pmos_5p04310591302027_3v256x8m81_2/S_uq0
+ pmos_5p04310591302027_3v256x8m81_2/S pmos_5p04310591302027_3v256x8m81
Xnmos_5p04310591302032_3v256x8m81_0 nmos_5p04310591302032_3v256x8m81_0/D nmos_5p04310591302034_3v256x8m81_0/D
+ nmos_5p04310591302034_3v256x8m81_0/D vss vss vss nmos_5p04310591302032_3v256x8m81
Xpmos_1p2$$46283820_3v256x8m81_0 pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ pcb pcb pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S pcb
+ pcb pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S vdd pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ vdd pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ vdd vdd pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S vdd
+ vdd vdd pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S pcb
+ pmos_1p2$$46283820_3v256x8m81
Xnmos_1p2$$45101100_3v256x8m81_0 men vss men vss vss men pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ men pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ men vss nmos_1p2$$45101100_3v256x8m81
Xnmos_5p04310591302033_3v256x8m81_0 vss pmos_5p04310591302027_3v256x8m81_0/S_uq0 pmos_5p04310591302038_3v256x8m81_0/S
+ vss nmos_5p04310591302033_3v256x8m81
Xpmos_1p2$$46287916_3v256x8m81_0 vdd vdd nmos_5p04310591302034_3v256x8m81_0/D nmos_5p04310591302032_3v256x8m81_0/D
+ vdd nmos_5p04310591302034_3v256x8m81_0/D pmos_1p2$$46287916_3v256x8m81
Xnmos_5p04310591302034_3v256x8m81_0 nmos_5p04310591302034_3v256x8m81_0/D pmos_5p04310591302027_3v256x8m81_1/S
+ vss vss nmos_5p04310591302034_3v256x8m81
Xpmos_1p2$$46284844_3v256x8m81_0 vdd_uq0 vdd_uq0 vdd_uq0 nmos_5p04310591302034_3v256x8m81_0/D
+ pmos_5p04310591302027_3v256x8m81_1/S pmos_5p04310591302027_3v256x8m81_1/S pmos_1p2$$46284844_3v256x8m81
Xnmos_1p2$$45102124_3v256x8m81_0 pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ vss pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S vss vss
+ vss pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S pcb pcb pcb
+ pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ pcb vss nmos_1p2$$45102124_3v256x8m81
Xpmos_1p2$$46286892_3v256x8m81_0 vdd vdd nmos_5p04310591302028_3v256x8m81_1/S nmos_5p04310591302028_3v256x8m81_1/S
+ nmos_5p04310591302032_3v256x8m81_0/D nmos_5p04310591302032_3v256x8m81_0/D nmos_5p04310591302032_3v256x8m81_0/D
+ vdd pmos_1p2$$46286892_3v256x8m81
Xnmos_5p04310591302023_3v256x8m81_0 vss pmos_5p04310591302027_3v256x8m81_2/S_uq0 pmos_5p04310591302027_3v256x8m81_0/S
+ pmos_5p04310591302027_3v256x8m81_0/S_uq0 pmos_5p04310591302027_3v256x8m81_0/S vss
+ nmos_5p04310591302023_3v256x8m81
Xnmos_5p04310591302028_3v256x8m81_0 nmos_5p04310591302028_3v256x8m81_1/D nmos_5p04310591302028_3v256x8m81_1/D
+ nmos_5p04310591302028_3v256x8m81_1/D nmos_5p04310591302032_3v256x8m81_0/D nmos_5p04310591302032_3v256x8m81_0/D
+ nmos_5p04310591302032_3v256x8m81_0/D nmos_5p04310591302032_3v256x8m81_0/D vss vss
+ vss nmos_5p04310591302032_3v256x8m81_0/D vss nmos_5p04310591302028_3v256x8m81
Xpmos_1p2$$46281772_3v256x8m81_0 pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S
+ pmos_1p2$$46281772_3v256x8m81_0/pmos_5p04310591302025_3v256x8m81_0/S pmos_1p2$$46281772_3v256x8m81_1/pmos_5p04310591302025_3v256x8m81_0/S
+ vdd pmos_1p2$$46281772_3v256x8m81_1/pmos_5p04310591302025_3v256x8m81_0/S vdd vdd
+ pmos_1p2$$46281772_3v256x8m81_1/pmos_5p04310591302025_3v256x8m81_0/S pmos_1p2$$46281772_3v256x8m81
Xnmos_5p04310591302023_3v256x8m81_1 vss pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ vss pmos_5p04310591302027_3v256x8m81_1/S_uq0 pmos_5p04310591302027_3v256x8m81_1/S
+ vss nmos_5p04310591302023_3v256x8m81
Xnmos_5p04310591302028_3v256x8m81_1 nmos_5p04310591302028_3v256x8m81_1/D nmos_5p04310591302028_3v256x8m81_1/D
+ nmos_5p04310591302028_3v256x8m81_1/D pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D nmos_5p04310591302028_3v256x8m81_1/S
+ nmos_5p04310591302028_3v256x8m81_1/S nmos_5p04310591302028_3v256x8m81_1/S pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ vss nmos_5p04310591302028_3v256x8m81
Xpmos_1p2$$46281772_3v256x8m81_1 pmos_1p2$$46281772_3v256x8m81_1/pmos_5p04310591302025_3v256x8m81_0/S
+ pmos_1p2$$46281772_3v256x8m81_1/pmos_5p04310591302025_3v256x8m81_0/S nmos_5p04310591302028_3v256x8m81_1/S
+ vdd pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D vdd vdd
+ nmos_5p04310591302034_3v256x8m81_0/D pmos_1p2$$46281772_3v256x8m81
Xnmos_5p04310591302023_3v256x8m81_2 vss pmos_5p04310591302027_3v256x8m81_1/S_uq0 pmos_5p04310591302027_3v256x8m81_2/S
+ pmos_5p04310591302027_3v256x8m81_2/S_uq0 pmos_5p04310591302027_3v256x8m81_2/S vss
+ nmos_5p04310591302023_3v256x8m81
Xpmos_1p2$$46285868_3v256x8m81_0 vdd nmos_5p04310591302028_3v256x8m81_1/S vdd pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ pmos_1p2$$46285868_3v256x8m81
Xpmos_5p04310591302038_3v256x8m81_0 vdd_uq0 pmos_5p04310591302027_3v256x8m81_0/S_uq0
+ vdd_uq0 pmos_5p04310591302038_3v256x8m81_0/S pmos_5p04310591302038_3v256x8m81
Xnmos_1p2$$45103148_3v256x8m81_0 nmos_5p04310591302028_3v256x8m81_1/S pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D
+ nmos_5p04310591302034_3v256x8m81_0/D vss vss nmos_5p04310591302028_3v256x8m81_1/S
+ nmos_5p04310591302034_3v256x8m81_0/D pmos_1p2$$46281772_3v256x8m81_1/pmos_5p04310591302025_3v256x8m81_0/S
+ pmos_1p2$$46282796_3v256x8m81_0/pmos_5p04310591302024_3v256x8m81_0/D vss nmos_1p2$$45103148_3v256x8m81
Xnmos_5p04310591302012_3v256x8m81_0 nmos_5p04310591302028_3v256x8m81_1/S se se nmos_5p04310591302028_3v256x8m81_1/S
+ vss vss vss nmos_5p04310591302028_3v256x8m81_1/S nmos_5p04310591302028_3v256x8m81_1/S
+ vss nmos_5p04310591302012_3v256x8m81
.ends

.subckt nmos_5p04310591302050_3v256x8m81 D_uq0 D a_265_n44# S_uq0 S a_n56_n44# a_104_n44#
+ VSUBS
X0 D_uq0 a_265_n44# S_uq0 VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.27692p ps=1.58u w=1.055u l=0.28u
X1 D a_n56_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X2 S_uq0 a_104_n44# D VSUBS nfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt nmos_5p04310591302044_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.451p pd=2.93u as=0.451p ps=2.93u w=1.025u l=0.28u
.ends

.subckt pmos_5p04310591302047_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.8206p pd=4.61u as=0.8206p ps=4.61u w=1.865u l=0.28u
.ends

.subckt nmos_5p0431059130208_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
.ends

.subckt nmos_5p04310591302045_3v256x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.583p ps=3.53u w=1.325u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.583p pd=3.53u as=0.3445p ps=1.845u w=1.325u l=0.28u
.ends

.subckt nmos_5p04310591302052_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.3278p pd=2.37u as=0.3278p ps=2.37u w=0.745u l=0.28u
.ends

.subckt pmos_5p04310591302048_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.924p pd=5.08u as=0.924p ps=5.08u w=2.1u l=0.28u
.ends

.subckt nmos_5p04310591302046_3v256x8m81 a_20_n44# D_uq1 D_uq0 D a_181_n44# a_502_n44#
+ S_uq2 a_662_n44# S_uq1 a_n140_n44# S_uq0 S a_341_n44# VSUBS
X0 S a_341_n44# D VSUBS nfet_03v3 ad=0.25855p pd=1.51u as=0.2561p ps=1.505u w=0.985u l=0.28u
X1 S_uq0 a_662_n44# D_uq0 VSUBS nfet_03v3 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.28u
X2 D_uq0 a_502_n44# S VSUBS nfet_03v3 ad=0.2561p pd=1.505u as=0.25855p ps=1.51u w=0.985u l=0.28u
X3 S_uq1 a_20_n44# D_uq1 VSUBS nfet_03v3 ad=0.25855p pd=1.51u as=0.2561p ps=1.505u w=0.985u l=0.28u
X4 D a_181_n44# S_uq1 VSUBS nfet_03v3 ad=0.2561p pd=1.505u as=0.25855p ps=1.51u w=0.985u l=0.28u
X5 D_uq1 a_n140_n44# S_uq2 VSUBS nfet_03v3 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.28u
.ends

.subckt pmos_5p04310591302049_3v256x8m81 a_20_n44# D_uq1 D_uq0 D a_181_n44# S_uq2
+ S_uq1 a_n140_n44# S_uq0 S a_341_n44# a_503_n44# a_663_n44# w_n314_n86#
X0 S a_341_n44# D w_n314_n86# pfet_03v3 ad=0.4664p pd=2.29u as=0.4576p ps=2.28u w=1.76u l=0.28u
X1 S_uq1 a_20_n44# D_uq1 w_n314_n86# pfet_03v3 ad=0.462p pd=2.285u as=0.4576p ps=2.28u w=1.76u l=0.28u
X2 D a_181_n44# S_uq1 w_n314_n86# pfet_03v3 ad=0.4576p pd=2.28u as=0.462p ps=2.285u w=1.76u l=0.28u
X3 D_uq1 a_n140_n44# S_uq2 w_n314_n86# pfet_03v3 ad=0.4576p pd=2.28u as=0.7744p ps=4.4u w=1.76u l=0.28u
X4 S_uq0 a_663_n44# D_uq0 w_n314_n86# pfet_03v3 ad=0.7832p pd=4.41u as=0.4576p ps=2.28u w=1.76u l=0.28u
X5 D_uq0 a_503_n44# S w_n314_n86# pfet_03v3 ad=0.4576p pd=2.28u as=0.4664p ps=2.29u w=1.76u l=0.28u
.ends

.subckt pmos_5p04310591302051_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.6877p pd=3.165u as=1.1638p ps=6.17u w=2.645u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=1.1638p pd=6.17u as=0.6877p ps=3.165u w=2.645u l=0.28u
.ends

.subckt pmos_5p0431059130203_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.1378p pd=1.05u as=0.2332p ps=1.94u w=0.53u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.2332p pd=1.94u as=0.1378p ps=1.05u w=0.53u l=0.28u
.ends

.subckt pmos_1p2$$171625516_3v256x8m81 a_n42_n34# pmos_5p0431059130203_3v256x8m81_0/S_uq0
+ pmos_5p0431059130203_3v256x8m81_0/S pmos_5p0431059130203_3v256x8m81_0/w_n202_n86#
+ a_118_n34# pmos_5p0431059130203_3v256x8m81_0/D
Xpmos_5p0431059130203_3v256x8m81_0 pmos_5p0431059130203_3v256x8m81_0/D a_n42_n34#
+ a_118_n34# pmos_5p0431059130203_3v256x8m81_0/w_n202_n86# pmos_5p0431059130203_3v256x8m81_0/S_uq0
+ pmos_5p0431059130203_3v256x8m81_0/S pmos_5p0431059130203_3v256x8m81
.ends

.subckt outbuf_oe_3v256x8m81 qp qn se q GWE vdd vss
Xnmos_5p04310591302050_3v256x8m81_0 nmos_5p0431059130208_3v256x8m81_1/S nmos_5p0431059130208_3v256x8m81_1/S
+ nmos_5p0431059130208_3v256x8m81_0/D pmos_5p04310591302051_3v256x8m81_0/D pmos_5p04310591302051_3v256x8m81_0/D
+ nmos_5p0431059130208_3v256x8m81_0/D nmos_5p0431059130208_3v256x8m81_0/D vss nmos_5p04310591302050_3v256x8m81
Xnmos_5p04310591302044_3v256x8m81_0 vss pmos_5p04310591302047_3v256x8m81_0/S pmos_5p04310591302048_3v256x8m81_0/S
+ vss nmos_5p04310591302044_3v256x8m81
Xpmos_5p04310591302047_3v256x8m81_0 vdd GWE vdd pmos_5p04310591302047_3v256x8m81_0/S
+ pmos_5p04310591302047_3v256x8m81
Xnmos_5p0431059130208_3v256x8m81_0 nmos_5p0431059130208_3v256x8m81_0/D se vss vss
+ nmos_5p0431059130208_3v256x8m81
Xnmos_5p0431059130208_3v256x8m81_1 vss pmos_5p04310591302038_3v256x8m81_0/D nmos_5p0431059130208_3v256x8m81_1/S
+ vss nmos_5p0431059130208_3v256x8m81
Xnmos_5p04310591302033_3v256x8m81_0 pmos_5p04310591302038_3v256x8m81_0/D pmos_5p04310591302051_3v256x8m81_0/D
+ vss vss nmos_5p04310591302033_3v256x8m81
Xnmos_5p04310591302045_3v256x8m81_0 vss pmos_5p04310591302047_3v256x8m81_0/S pmos_5p04310591302047_3v256x8m81_0/S
+ nmos_5p04310591302045_3v256x8m81_1/S nmos_5p04310591302045_3v256x8m81_1/S vss nmos_5p04310591302045_3v256x8m81
Xnmos_5p04310591302045_3v256x8m81_1 pmos_5p04310591302051_3v256x8m81_0/D qn qn nmos_5p04310591302045_3v256x8m81_1/S
+ nmos_5p04310591302045_3v256x8m81_1/S vss nmos_5p04310591302045_3v256x8m81
Xnmos_5p04310591302052_3v256x8m81_0 vss GWE pmos_5p04310591302047_3v256x8m81_0/S vss
+ nmos_5p04310591302052_3v256x8m81
Xpmos_5p04310591302048_3v256x8m81_0 vdd pmos_5p04310591302047_3v256x8m81_0/S vdd pmos_5p04310591302048_3v256x8m81_0/S
+ pmos_5p04310591302048_3v256x8m81
Xpmos_5p04310591302013_3v256x8m81_0 nmos_5p0431059130208_3v256x8m81_1/S nmos_5p0431059130208_3v256x8m81_1/S
+ se pmos_5p04310591302051_3v256x8m81_0/D pmos_5p04310591302051_3v256x8m81_0/D se
+ se vdd pmos_5p04310591302013_3v256x8m81
Xnmos_5p04310591302046_3v256x8m81_0 pmos_5p04310591302051_3v256x8m81_0/D vss vss vss
+ pmos_5p04310591302051_3v256x8m81_0/D pmos_5p04310591302051_3v256x8m81_0/D q pmos_5p04310591302051_3v256x8m81_0/D
+ q pmos_5p04310591302051_3v256x8m81_0/D q q pmos_5p04310591302051_3v256x8m81_0/D
+ vss nmos_5p04310591302046_3v256x8m81
Xpmos_5p04310591302049_3v256x8m81_0 pmos_5p04310591302051_3v256x8m81_0/D vdd vdd vdd
+ pmos_5p04310591302051_3v256x8m81_0/D q q pmos_5p04310591302051_3v256x8m81_0/D q
+ q pmos_5p04310591302051_3v256x8m81_0/D pmos_5p04310591302051_3v256x8m81_0/D pmos_5p04310591302051_3v256x8m81_0/D
+ vdd pmos_5p04310591302049_3v256x8m81
Xpmos_5p04310591302051_3v256x8m81_0 pmos_5p04310591302051_3v256x8m81_0/D qp qp vdd
+ pmos_5p04310591302051_3v256x8m81_1/S pmos_5p04310591302051_3v256x8m81_1/S pmos_5p04310591302051_3v256x8m81
Xpmos_5p04310591302051_3v256x8m81_1 vdd pmos_5p04310591302048_3v256x8m81_0/S pmos_5p04310591302048_3v256x8m81_0/S
+ vdd pmos_5p04310591302051_3v256x8m81_1/S pmos_5p04310591302051_3v256x8m81_1/S pmos_5p04310591302051_3v256x8m81
Xpmos_1p2$$171625516_3v256x8m81_0 pmos_5p04310591302038_3v256x8m81_0/D vdd vdd vdd
+ pmos_5p04310591302038_3v256x8m81_0/D nmos_5p0431059130208_3v256x8m81_1/S pmos_1p2$$171625516_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_0 nmos_5p0431059130208_3v256x8m81_0/D se vdd vdd
+ pmos_5p04310591302014_3v256x8m81
Xpmos_5p04310591302038_3v256x8m81_0 pmos_5p04310591302038_3v256x8m81_0/D pmos_5p04310591302051_3v256x8m81_0/D
+ vdd vdd pmos_5p04310591302038_3v256x8m81
.ends

.subckt pmos_5p0431059130209_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.3276p pd=11.46u as=2.3276p ps=11.46u w=5.29u l=0.28u
.ends

.subckt nmos_5p0431059130207_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=2.794p pd=13.58u as=2.794p ps=13.58u w=6.35u l=0.28u
.ends

.subckt nmos_1p2$$46884908_3v256x8m81 nmos_5p0431059130207_3v256x8m81_0/S a_n14_n34#
+ nmos_5p0431059130207_3v256x8m81_0/D VSUBS
Xnmos_5p0431059130207_3v256x8m81_0 nmos_5p0431059130207_3v256x8m81_0/D a_n14_n34#
+ nmos_5p0431059130207_3v256x8m81_0/S VSUBS nmos_5p0431059130207_3v256x8m81
.ends

.subckt pmos_5p0431059130201_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=1.397p pd=7.23u as=1.397p ps=7.23u w=3.175u l=0.28u
.ends

.subckt pmos_1p2$$46889004_3v256x8m81 pmos_5p0431059130201_3v256x8m81_0/D a_n14_n34#
+ pmos_5p0431059130201_3v256x8m81_0/S w_n133_n66#
Xpmos_5p0431059130201_3v256x8m81_0 pmos_5p0431059130201_3v256x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p0431059130201_3v256x8m81_0/S pmos_5p0431059130201_3v256x8m81
.ends

.subckt nmos_5p0431059130205_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=2.3276p pd=11.46u as=2.3276p ps=11.46u w=5.29u l=0.28u
.ends

.subckt nmos_1p2$$46883884_3v256x8m81 nmos_5p0431059130205_3v256x8m81_0/D a_n14_n34#
+ nmos_5p0431059130205_3v256x8m81_0/S VSUBS
Xnmos_5p0431059130205_3v256x8m81_0 nmos_5p0431059130205_3v256x8m81_0/D a_n14_n34#
+ nmos_5p0431059130205_3v256x8m81_0/S VSUBS nmos_5p0431059130205_3v256x8m81
.ends

.subckt pmos_5p0431059130206_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.1157p pd=0.965u as=0.1958p ps=1.77u w=0.445u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.1958p pd=1.77u as=0.1157p ps=0.965u w=0.445u l=0.28u
.ends

.subckt nmos_5p04310591302010_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.4642p ps=2.99u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46273580_3v256x8m81 w_n133_n66# a_n42_n34# pmos_5p0431059130203_3v256x8m81_0/S
+ pmos_5p0431059130203_3v256x8m81_0/S_uq0 a_118_n34# pmos_5p0431059130203_3v256x8m81_0/D
Xpmos_5p0431059130203_3v256x8m81_0 pmos_5p0431059130203_3v256x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p0431059130203_3v256x8m81_0/S_uq0 pmos_5p0431059130203_3v256x8m81_0/S
+ pmos_5p0431059130203_3v256x8m81
.ends

.subckt nmos_5p04310591302011_3v256x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.1157p pd=0.965u as=0.1958p ps=1.77u w=0.445u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.1958p pd=1.77u as=0.1157p ps=0.965u w=0.445u l=0.28u
.ends

.subckt pmos_1p2$$46885932_3v256x8m81 pmos_5p0431059130206_3v256x8m81_0/S pmos_5p0431059130206_3v256x8m81_0/D
+ pmos_5p0431059130206_3v256x8m81_0/S_uq0 a_118_89# a_n42_89# w_n133_n65#
Xpmos_5p0431059130206_3v256x8m81_0 pmos_5p0431059130206_3v256x8m81_0/D a_n42_89# a_118_89#
+ w_n133_n65# pmos_5p0431059130206_3v256x8m81_0/S_uq0 pmos_5p0431059130206_3v256x8m81_0/S
+ pmos_5p0431059130206_3v256x8m81
.ends

.subckt nmos_1p2$$46563372_3v256x8m81 nmos_5p0431059130208_3v256x8m81_0/D a_n14_89#
+ nmos_5p0431059130208_3v256x8m81_0/S VSUBS
Xnmos_5p0431059130208_3v256x8m81_0 nmos_5p0431059130208_3v256x8m81_0/D a_n14_89# nmos_5p0431059130208_3v256x8m81_0/S
+ VSUBS nmos_5p0431059130208_3v256x8m81
.ends

.subckt pmos_5p0431059130204_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.794p pd=13.58u as=2.794p ps=13.58u w=6.35u l=0.28u
.ends

.subckt pmos_1p2$$46887980_3v256x8m81 w_n133_n66# pmos_5p0431059130204_3v256x8m81_0/S
+ a_n14_n34# pmos_5p0431059130204_3v256x8m81_0/D
Xpmos_5p0431059130204_3v256x8m81_0 pmos_5p0431059130204_3v256x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p0431059130204_3v256x8m81_0/S pmos_5p0431059130204_3v256x8m81
.ends

.subckt din_3v256x8m81 vss datain men db d wep vdd pmos_5p0431059130206_3v256x8m81_0/D
+ m1_114_5647# VSUBS
Xpmos_5p0431059130209_3v256x8m81_0 vdd pmos_1p2$$46889004_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ vdd pmos_5p0431059130209_3v256x8m81_0/S pmos_5p0431059130209_3v256x8m81
Xnmos_1p2$$46884908_3v256x8m81_0 VSUBS pmos_5p0431059130201_3v256x8m81_0/S pmos_1p2$$46889004_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ VSUBS nmos_1p2$$46884908_3v256x8m81
Xpmos_1p2$$46889004_3v256x8m81_0 pmos_1p2$$46889004_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ a_507_5030# d vdd pmos_1p2$$46889004_3v256x8m81
Xpmos_5p0431059130201_3v256x8m81_0 pmos_5p0431059130206_3v256x8m81_0/D nmos_5p04310591302011_3v256x8m81_1/D
+ pmos_5p0431059130206_3v256x8m81_0/D pmos_5p0431059130201_3v256x8m81_0/S pmos_5p0431059130201_3v256x8m81
Xnmos_1p2$$46883884_3v256x8m81_0 pmos_5p0431059130209_3v256x8m81_0/S wep db VSUBS
+ nmos_1p2$$46883884_3v256x8m81
Xpmos_1p2$$46889004_3v256x8m81_1 pmos_5p0431059130209_3v256x8m81_0/S a_507_5030# db
+ vdd pmos_1p2$$46889004_3v256x8m81
Xpmos_5p0431059130206_3v256x8m81_0 pmos_5p0431059130206_3v256x8m81_0/D datain pmos_5p0431059130206_3v256x8m81_0/S
+ pmos_5p0431059130206_3v256x8m81_0/D nmos_5p04310591302011_3v256x8m81_1/S pmos_5p0431059130206_3v256x8m81_0/S
+ pmos_5p0431059130206_3v256x8m81
Xnmos_1p2$$46883884_3v256x8m81_1 VSUBS pmos_1p2$$46889004_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ pmos_5p0431059130209_3v256x8m81_0/S VSUBS nmos_1p2$$46883884_3v256x8m81
Xnmos_5p04310591302010_3v256x8m81_0 VSUBS nmos_5p04310591302011_3v256x8m81_1/D pmos_5p0431059130201_3v256x8m81_0/S
+ VSUBS nmos_5p04310591302010_3v256x8m81
Xpmos_1p2$$46273580_3v256x8m81_0 pmos_5p0431059130206_3v256x8m81_0/D men pmos_5p0431059130206_3v256x8m81_0/D
+ pmos_5p0431059130206_3v256x8m81_0/D men pmos_1p2$$46273580_3v256x8m81_0/pmos_5p0431059130203_3v256x8m81_0/D
+ pmos_1p2$$46273580_3v256x8m81
Xnmos_1p2$$46883884_3v256x8m81_2 pmos_1p2$$46889004_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ wep d VSUBS nmos_1p2$$46883884_3v256x8m81
Xpmos_1p2$$46273580_3v256x8m81_1 pmos_5p0431059130206_3v256x8m81_0/D pmos_5p0431059130201_3v256x8m81_0/S
+ pmos_5p0431059130206_3v256x8m81_0/D pmos_5p0431059130206_3v256x8m81_0/D pmos_5p0431059130201_3v256x8m81_0/S
+ nmos_5p04310591302011_3v256x8m81_1/S_uq0 pmos_1p2$$46273580_3v256x8m81
Xnmos_5p04310591302011_3v256x8m81_0 VSUBS datain pmos_5p0431059130206_3v256x8m81_0/S
+ nmos_5p04310591302011_3v256x8m81_1/S pmos_5p0431059130206_3v256x8m81_0/S VSUBS nmos_5p04310591302011_3v256x8m81
Xnmos_5p04310591302011_3v256x8m81_1 nmos_5p04310591302011_3v256x8m81_1/D pmos_1p2$$46273580_3v256x8m81_0/pmos_5p0431059130203_3v256x8m81_0/D
+ men nmos_5p04310591302011_3v256x8m81_1/S_uq0 nmos_5p04310591302011_3v256x8m81_1/S
+ VSUBS nmos_5p04310591302011_3v256x8m81
Xpmos_1p2$$46885932_3v256x8m81_0 nmos_5p04310591302011_3v256x8m81_1/S nmos_5p04310591302011_3v256x8m81_1/D
+ nmos_5p04310591302011_3v256x8m81_1/S_uq0 pmos_1p2$$46273580_3v256x8m81_0/pmos_5p0431059130203_3v256x8m81_0/D
+ men pmos_5p0431059130206_3v256x8m81_0/D pmos_1p2$$46885932_3v256x8m81
Xnmos_1p2$$46563372_3v256x8m81_0 nmos_5p04310591302011_3v256x8m81_1/S_uq0 pmos_5p0431059130201_3v256x8m81_0/S
+ VSUBS VSUBS nmos_1p2$$46563372_3v256x8m81
Xnmos_1p2$$46563372_3v256x8m81_1 pmos_1p2$$46273580_3v256x8m81_0/pmos_5p0431059130203_3v256x8m81_0/D
+ men VSUBS VSUBS nmos_1p2$$46563372_3v256x8m81
Xpmos_1p2$$46887980_3v256x8m81_0 vdd vdd pmos_5p0431059130201_3v256x8m81_0/S pmos_1p2$$46889004_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ pmos_1p2$$46887980_3v256x8m81
X0 vdd wep a_507_5030# vdd pfet_03v3 ad=0.38572p pd=2.5u as=0.1859p ps=1.23u w=0.695u l=0.28u
X1 a_507_5030# wep vdd vdd pfet_03v3 ad=0.1859p pd=1.23u as=0.38572p ps=2.5u w=0.695u l=0.28u
X2 a_507_5030# wep vss VSUBS nfet_03v3 ad=0.28355p pd=2.13u as=0.3103p ps=2.23u w=0.535u l=0.28u
.ends

.subckt nmos_1p2$$202596396_3v256x8m81 nmos_5p0431059130208_3v256x8m81_0/D a_n14_89#
+ nmos_5p0431059130208_3v256x8m81_0/S VSUBS
Xnmos_5p0431059130208_3v256x8m81_0 nmos_5p0431059130208_3v256x8m81_0/D a_n14_89# nmos_5p0431059130208_3v256x8m81_0/S
+ VSUBS nmos_5p0431059130208_3v256x8m81
.ends

.subckt pmos_5p04310591302041_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.1958p pd=1.77u as=0.1958p ps=1.77u w=0.445u l=0.28u
.ends

.subckt nmos_5p04310591302040_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.2794p pd=2.15u as=0.2794p ps=2.15u w=0.635u l=0.28u
.ends

.subckt pmos_1p2$$202585132_3v256x8m81 pmos_5p04310591302014_3v256x8m81_0/S a_n14_n34#
+ pmos_5p04310591302014_3v256x8m81_0/D w_n119_n65#
Xpmos_5p04310591302014_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_0/D a_n14_n34#
+ w_n119_n65# pmos_5p04310591302014_3v256x8m81_0/S pmos_5p04310591302014_3v256x8m81
.ends

.subckt pmos_5p04310591302043_3v256x8m81 D_uq0 D a_265_n44# S_uq0 S a_n56_n44# a_104_n44#
+ w_n230_n86#
X0 D_uq0 a_265_n44# S_uq0 w_n230_n86# pfet_03v3 ad=0.4092p pd=2.74u as=0.24412p ps=1.455u w=0.93u l=0.28u
X1 D a_n56_n44# S w_n230_n86# pfet_03v3 ad=0.2418p pd=1.45u as=0.4092p ps=2.74u w=0.93u l=0.28u
X2 S_uq0 a_104_n44# D w_n230_n86# pfet_03v3 ad=0.24412p pd=1.455u as=0.2418p ps=1.45u w=0.93u l=0.28u
.ends

.subckt nmos_1p2$$202598444_3v256x8m81 nmos_5p04310591302010_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v256x8m81_0/S VSUBS
Xnmos_5p04310591302010_3v256x8m81_0 nmos_5p04310591302010_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v256x8m81_0/S VSUBS nmos_5p04310591302010_3v256x8m81
.ends

.subckt pmos_1p2$$202587180_3v256x8m81 pmos_5p04310591302014_3v256x8m81_0/S a_n14_n34#
+ pmos_5p04310591302014_3v256x8m81_0/D w_n133_n65#
Xpmos_5p04310591302014_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302014_3v256x8m81_0/S pmos_5p04310591302014_3v256x8m81
.ends

.subckt pmos_1p2$$202584108_3v256x8m81 pmos_5p04310591302014_3v256x8m81_0/S a_n14_n34#
+ pmos_5p04310591302014_3v256x8m81_0/D w_n133_n65#
Xpmos_5p04310591302014_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302014_3v256x8m81_0/S pmos_5p04310591302014_3v256x8m81
.ends

.subckt pmos_5p04310591302020_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt nmos_5p04310591302039_3v256x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.4642p pd=2.99u as=0.2743p ps=1.575u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$202586156_3v256x8m81 pmos_5p04310591302014_3v256x8m81_0/S a_n14_n34#
+ pmos_5p04310591302014_3v256x8m81_0/D w_n133_n65#
Xpmos_5p04310591302014_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302014_3v256x8m81_0/S pmos_5p04310591302014_3v256x8m81
.ends

.subckt nmos_1p2$$202595372_3v256x8m81 nmos_5p0431059130208_3v256x8m81_0/D a_n14_89#
+ nmos_5p0431059130208_3v256x8m81_0/S VSUBS
Xnmos_5p0431059130208_3v256x8m81_0 nmos_5p0431059130208_3v256x8m81_0/D a_n14_89# nmos_5p0431059130208_3v256x8m81_0/S
+ VSUBS nmos_5p0431059130208_3v256x8m81
.ends

.subckt nmos_5p04310591302042_3v256x8m81 D_uq0 D a_265_n44# S_uq0 S a_n56_n44# a_104_n44#
+ VSUBS
X0 D_uq0 a_265_n44# S_uq0 VSUBS nfet_03v3 ad=0.1628p pd=1.62u as=97.125f ps=0.895u w=0.37u l=0.28u
X1 D a_n56_n44# S VSUBS nfet_03v3 ad=96.2f pd=0.89u as=0.1628p ps=1.62u w=0.37u l=0.28u
X2 S_uq0 a_104_n44# D VSUBS nfet_03v3 ad=97.125f pd=0.895u as=96.2f ps=0.89u w=0.37u l=0.28u
.ends

.subckt nmos_1p2$$202594348_3v256x8m81 nmos_5p04310591302040_3v256x8m81_0/S nmos_5p04310591302040_3v256x8m81_0/D
+ a_n14_n44# VSUBS
Xnmos_5p04310591302040_3v256x8m81_0 nmos_5p04310591302040_3v256x8m81_0/D a_n14_n44#
+ nmos_5p04310591302040_3v256x8m81_0/S VSUBS nmos_5p04310591302040_3v256x8m81
.ends

.subckt pmos_1p2$$202583084_3v256x8m81 a_n42_n34# pmos_5p04310591302035_3v256x8m81_0/S
+ pmos_5p04310591302035_3v256x8m81_0/S_uq0 w_n133_n66# pmos_5p04310591302035_3v256x8m81_0/D
+ a_118_n34#
Xpmos_5p04310591302035_3v256x8m81_0 pmos_5p04310591302035_3v256x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302035_3v256x8m81_0/S_uq0 pmos_5p04310591302035_3v256x8m81_0/S
+ pmos_5p04310591302035_3v256x8m81
.ends

.subckt wen_wm1_3v256x8m81 GWEN men wep vss vdd wen vdd_uq0
Xnmos_1p2$$202596396_3v256x8m81_0 nmos_1p2$$202596396_3v256x8m81_0/nmos_5p0431059130208_3v256x8m81_0/D
+ nmos_1p2$$202595372_3v256x8m81_1/nmos_5p0431059130208_3v256x8m81_0/S vss vss nmos_1p2$$202596396_3v256x8m81
Xnmos_1p2$$202596396_3v256x8m81_1 vss nmos_1p2$$202595372_3v256x8m81_1/nmos_5p0431059130208_3v256x8m81_0/S
+ pmos_5p04310591302041_3v256x8m81_0/D vss nmos_1p2$$202596396_3v256x8m81
Xpmos_5p04310591302041_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_0/D pmos_5p04310591302014_3v256x8m81_5/D
+ vdd pmos_5p04310591302041_3v256x8m81_0/S pmos_5p04310591302041_3v256x8m81
Xpmos_5p04310591302035_3v256x8m81_0 pmos_5p04310591302035_3v256x8m81_0/D pmos_5p04310591302020_3v256x8m81_0/S
+ pmos_5p04310591302020_3v256x8m81_0/S vdd_uq0 vdd_uq0 vdd_uq0 pmos_5p04310591302035_3v256x8m81
Xnmos_5p0431059130208_3v256x8m81_0 vss GWEN nmos_5p0431059130208_3v256x8m81_2/D vss
+ nmos_5p0431059130208_3v256x8m81
Xnmos_5p0431059130208_3v256x8m81_1 nmos_5p0431059130208_3v256x8m81_1/D nmos_5p0431059130208_3v256x8m81_2/D
+ vss vss nmos_5p0431059130208_3v256x8m81
Xnmos_5p0431059130208_3v256x8m81_2 nmos_5p0431059130208_3v256x8m81_2/D wen vss vss
+ nmos_5p0431059130208_3v256x8m81
Xnmos_5p04310591302040_3v256x8m81_0 pmos_5p04310591302035_3v256x8m81_0/D pmos_5p04310591302020_3v256x8m81_0/S
+ vss vss nmos_5p04310591302040_3v256x8m81
Xnmos_5p0431059130208_3v256x8m81_3 nmos_5p0431059130208_3v256x8m81_3/D pmos_5p04310591302014_3v256x8m81_5/D
+ vss vss nmos_5p0431059130208_3v256x8m81
Xnmos_5p04310591302040_3v256x8m81_1 pmos_5p04310591302014_3v256x8m81_5/D men vss vss
+ nmos_5p04310591302040_3v256x8m81
Xpmos_1p2$$202585132_3v256x8m81_0 vdd nmos_1p2$$202595372_3v256x8m81_1/nmos_5p0431059130208_3v256x8m81_0/S
+ nmos_1p2$$202596396_3v256x8m81_0/nmos_5p0431059130208_3v256x8m81_0/D vdd pmos_1p2$$202585132_3v256x8m81
Xnmos_5p04310591302040_3v256x8m81_2 vss vss pmos_5p04310591302014_3v256x8m81_5/D vss
+ nmos_5p04310591302040_3v256x8m81
Xpmos_5p04310591302043_3v256x8m81_0 wep wep pmos_5p04310591302035_3v256x8m81_0/D vdd_uq0
+ vdd_uq0 pmos_5p04310591302035_3v256x8m81_0/D pmos_5p04310591302035_3v256x8m81_0/D
+ vdd_uq0 pmos_5p04310591302043_3v256x8m81
Xnmos_5p04310591302010_3v256x8m81_0 vss nmos_1p2$$202596396_3v256x8m81_0/nmos_5p0431059130208_3v256x8m81_0/D
+ pmos_5p04310591302020_3v256x8m81_0/S vss nmos_5p04310591302010_3v256x8m81
Xnmos_1p2$$202598444_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_0/S pmos_5p04310591302014_3v256x8m81_5/D
+ nmos_5p0431059130208_3v256x8m81_1/D vss nmos_1p2$$202598444_3v256x8m81
Xpmos_1p2$$202587180_3v256x8m81_0 nmos_5p0431059130208_3v256x8m81_1/D nmos_5p0431059130208_3v256x8m81_3/D
+ pmos_5p04310591302041_3v256x8m81_0/S vdd pmos_1p2$$202587180_3v256x8m81
Xpmos_1p2$$202584108_3v256x8m81_0 nmos_1p2$$202595372_3v256x8m81_1/nmos_5p0431059130208_3v256x8m81_0/S
+ pmos_5p04310591302041_3v256x8m81_0/S vdd vdd pmos_1p2$$202584108_3v256x8m81
Xpmos_5p04310591302020_3v256x8m81_0 men nmos_1p2$$202596396_3v256x8m81_0/nmos_5p0431059130208_3v256x8m81_0/D
+ nmos_1p2$$202596396_3v256x8m81_0/nmos_5p0431059130208_3v256x8m81_0/D vdd pmos_5p04310591302020_3v256x8m81_0/S
+ pmos_5p04310591302020_3v256x8m81_0/S pmos_5p04310591302020_3v256x8m81
Xnmos_5p04310591302039_3v256x8m81_0 men pmos_1p2$$202583084_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D
+ pmos_1p2$$202583084_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D pmos_5p04310591302020_3v256x8m81_0/S
+ pmos_5p04310591302020_3v256x8m81_0/S vss nmos_5p04310591302039_3v256x8m81
Xpmos_1p2$$202586156_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_0/D nmos_1p2$$202595372_3v256x8m81_1/nmos_5p0431059130208_3v256x8m81_0/S
+ vdd vdd pmos_1p2$$202586156_3v256x8m81
Xnmos_1p2$$202595372_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_0/D nmos_5p0431059130208_3v256x8m81_3/D
+ pmos_5p04310591302041_3v256x8m81_0/S vss nmos_1p2$$202595372_3v256x8m81
Xnmos_1p2$$202595372_3v256x8m81_1 vss pmos_5p04310591302041_3v256x8m81_0/S nmos_1p2$$202595372_3v256x8m81_1/nmos_5p0431059130208_3v256x8m81_0/S
+ vss nmos_1p2$$202595372_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_2/S wen vdd_uq0
+ vdd_uq0 pmos_5p04310591302014_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_1 nmos_5p0431059130208_3v256x8m81_1/D nmos_5p0431059130208_3v256x8m81_2/D
+ vdd_uq0 vdd_uq0 pmos_5p04310591302014_3v256x8m81
Xnmos_5p04310591302042_3v256x8m81_0 wep wep pmos_5p04310591302035_3v256x8m81_0/D vss
+ vss pmos_5p04310591302035_3v256x8m81_0/D pmos_5p04310591302035_3v256x8m81_0/D vss
+ nmos_5p04310591302042_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_2 nmos_5p0431059130208_3v256x8m81_2/D GWEN vdd_uq0
+ pmos_5p04310591302014_3v256x8m81_2/S pmos_5p04310591302014_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_3 pmos_5p04310591302014_3v256x8m81_5/S men vdd vdd
+ pmos_5p04310591302014_3v256x8m81
Xnmos_1p2$$202594348_3v256x8m81_0 pmos_1p2$$202583084_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D
+ vss nmos_1p2$$202596396_3v256x8m81_0/nmos_5p0431059130208_3v256x8m81_0/D vss nmos_1p2$$202594348_3v256x8m81
Xpmos_1p2$$202583084_3v256x8m81_0 nmos_1p2$$202596396_3v256x8m81_0/nmos_5p0431059130208_3v256x8m81_0/D
+ vdd vdd vdd pmos_1p2$$202583084_3v256x8m81_0/pmos_5p04310591302035_3v256x8m81_0/D
+ nmos_1p2$$202596396_3v256x8m81_0/nmos_5p0431059130208_3v256x8m81_0/D pmos_1p2$$202583084_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_4 nmos_5p0431059130208_3v256x8m81_3/D pmos_5p04310591302014_3v256x8m81_5/D
+ vdd vdd pmos_5p04310591302014_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_5 pmos_5p04310591302014_3v256x8m81_5/D vss vdd pmos_5p04310591302014_3v256x8m81_5/S
+ pmos_5p04310591302014_3v256x8m81
.ends

.subckt nmos_5p0431059130200_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.397p pd=7.23u as=1.397p ps=7.23u w=3.175u l=0.28u
.ends

.subckt nmos_1p2$$47119404_3v256x8m81 nmos_5p0431059130200_3v256x8m81_0/D a_n14_n34#
+ nmos_5p0431059130200_3v256x8m81_0/S VSUBS
Xnmos_5p0431059130200_3v256x8m81_0 nmos_5p0431059130200_3v256x8m81_0/D a_n14_n34#
+ nmos_5p0431059130200_3v256x8m81_0/S VSUBS nmos_5p0431059130200_3v256x8m81
.ends

.subckt nmos_5p0431059130202_3v256x8m81 D a_n32_n44# a_136_n44# S_uq0 S VSUBS
X0 D a_n32_n44# S VSUBS nfet_03v3 ad=91.3f pd=0.92u as=0.1561p ps=1.64u w=0.265u l=0.28u
X1 S_uq0 a_136_n44# D VSUBS nfet_03v3 ad=0.15742p pd=1.65u as=91.3f ps=0.92u w=0.265u l=0.28u
.ends

.subckt ypass_gate_3v256x8m81 vss vdd b bb ypass pcb vdd_uq0 m3_n41_6881# m3_n41_5924#
+ m3_n41_6639# m3_n41_4610# pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ m3_n41_5682# m3_n41_5198# m3_n41_5440# m3_n41_6156# VSUBS db
Xnmos_1p2$$47119404_3v256x8m81_1 pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass b VSUBS nmos_1p2$$47119404_3v256x8m81
Xnmos_1p2$$47119404_3v256x8m81_3 db ypass bb VSUBS nmos_1p2$$47119404_3v256x8m81
Xnmos_5p0431059130202_3v256x8m81_0 nmos_5p0431059130202_3v256x8m81_0/D ypass ypass
+ VSUBS VSUBS VSUBS nmos_5p0431059130202_3v256x8m81
Xpmos_5p0431059130201_3v256x8m81_0 b pcb vdd bb pmos_5p0431059130201_3v256x8m81
Xpmos_1p2$$46889004_3v256x8m81_1 pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ nmos_5p0431059130202_3v256x8m81_0/D b vdd_uq0 pmos_1p2$$46889004_3v256x8m81
Xpmos_5p0431059130201_3v256x8m81_1 db nmos_5p0431059130202_3v256x8m81_0/D vdd bb pmos_5p0431059130201_3v256x8m81
X0 vdd pcb b vdd pfet_03v3 ad=0.92722p pd=4.34u as=0.4121p ps=2.105u w=1.585u l=0.28u
X1 b pcb vdd vdd pfet_03v3 ad=0.4121p pd=2.105u as=0.93515p ps=4.35u w=1.585u l=0.28u
X2 nmos_5p0431059130202_3v256x8m81_0/D ypass vdd_uq0 vdd_uq0 pfet_03v3 ad=0.26235p pd=1.45u as=0.46218p ps=2.72u w=0.695u l=0.28u
X3 vdd_uq0 ypass nmos_5p0431059130202_3v256x8m81_0/D vdd_uq0 pfet_03v3 ad=0.39963p pd=2.54u as=0.26235p ps=1.45u w=0.695u l=0.28u
X4 vdd pcb bb vdd pfet_03v3 ad=0.93015p pd=4.35u as=0.4134p ps=2.11u w=1.59u l=0.28u
X5 bb pcb vdd vdd pfet_03v3 ad=0.4134p pd=2.11u as=0.9381p ps=4.36u w=1.59u l=0.28u
.ends

.subckt ypass_gate_a_3v256x8m81 vss b bb ypass pcb vdd_uq0 m3_n41_6881# m3_n41_5924#
+ m3_n41_6639# m3_n41_4610# m3_n41_5682# vdd pmos_5p0431059130201_3v256x8m81_0/D VSUBS
+ pmos_5p0431059130201_3v256x8m81_1/D pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ m3_n41_5198# m3_n41_5440# m3_n41_6156#
Xnmos_1p2$$47119404_3v256x8m81_1 pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass pmos_5p0431059130201_3v256x8m81_0/D VSUBS nmos_1p2$$47119404_3v256x8m81
Xnmos_1p2$$47119404_3v256x8m81_3 pmos_5p0431059130201_3v256x8m81_1/D ypass bb VSUBS
+ nmos_1p2$$47119404_3v256x8m81
Xnmos_5p0431059130202_3v256x8m81_0 nmos_5p0431059130202_3v256x8m81_0/D ypass ypass
+ VSUBS VSUBS VSUBS nmos_5p0431059130202_3v256x8m81
Xpmos_5p0431059130201_3v256x8m81_0 pmos_5p0431059130201_3v256x8m81_0/D pcb vdd bb
+ pmos_5p0431059130201_3v256x8m81
Xpmos_1p2$$46889004_3v256x8m81_1 pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ nmos_5p0431059130202_3v256x8m81_0/D pmos_5p0431059130201_3v256x8m81_0/D vdd_uq0
+ pmos_1p2$$46889004_3v256x8m81
Xpmos_5p0431059130201_3v256x8m81_1 pmos_5p0431059130201_3v256x8m81_1/D nmos_5p0431059130202_3v256x8m81_0/D
+ vdd bb pmos_5p0431059130201_3v256x8m81
X0 vdd pcb pmos_5p0431059130201_3v256x8m81_0/D vdd pfet_03v3 ad=1.06988p pd=4.52u as=0.4121p ps=2.105u w=1.585u l=0.28u
X1 pmos_5p0431059130201_3v256x8m81_0/D pcb vdd vdd pfet_03v3 ad=0.4121p pd=2.105u as=0.99855p ps=4.43u w=1.585u l=0.28u
X2 vdd_uq0 ypass nmos_5p0431059130202_3v256x8m81_0/D vdd_uq0 pfet_03v3 ad=0.5143p pd=2.87u as=0.34055p ps=1.675u w=0.695u l=0.28u
X3 vdd pcb bb vdd pfet_03v3 ad=1.07325p pd=4.53u as=0.4134p ps=2.11u w=1.59u l=0.28u
X4 bb pcb vdd vdd pfet_03v3 ad=0.4134p pd=2.11u as=1.0017p ps=4.44u w=1.59u l=0.28u
X5 nmos_5p0431059130202_3v256x8m81_0/D ypass vdd_uq0 vdd_uq0 pfet_03v3 ad=0.34055p pd=1.675u as=0.38572p ps=2.5u w=0.695u l=0.28u
.ends

.subckt mux821_3v256x8m81 ypass_gate_3v256x8m81_6/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_6/b ypass_gate_a_3v256x8m81_0/ypass ypass_gate_3v256x8m81_7/bb
+ ypass_gate_3v256x8m81_4/bb ypass_gate_3v256x8m81_1/bb ypass_gate_3v256x8m81_1/b
+ ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D ypass_gate_3v256x8m81_1/db
+ ypass_gate_3v256x8m81_1/ypass ypass_gate_3v256x8m81_7/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_4/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_3/b ypass_gate_3v256x8m81_2/ypass ypass_gate_3v256x8m81_3/ypass
+ ypass_gate_3v256x8m81_4/ypass ypass_gate_3v256x8m81_5/b ypass_gate_3v256x8m81_5/ypass
+ ypass_gate_3v256x8m81_6/ypass ypass_gate_3v256x8m81_7/ypass ypass_gate_3v256x8m81_7/b
+ ypass_gate_3v256x8m81_6/bb ypass_gate_3v256x8m81_3/bb ypass_gate_3v256x8m81_7/db
+ ypass_gate_3v256x8m81_5/db ypass_gate_3v256x8m81_5/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_a_3v256x8m81_0/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_a_3v256x8m81_0/bb ypass_gate_3v256x8m81_2/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5924# ypass_gate_3v256x8m81_7/pcb
+ ypass_gate_3v256x8m81_7/vss ypass_gate_3v256x8m81_7/m3_n41_5440# ypass_gate_3v256x8m81_2/b
+ ypass_gate_3v256x8m81_7/vdd ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_7/m3_n41_6156#
+ ypass_gate_3v256x8m81_5/bb ypass_gate_3v256x8m81_2/bb ypass_gate_3v256x8m81_4/b
+ ypass_gate_3v256x8m81_3/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_1/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ VSUBS ypass_gate_3v256x8m81_4/db ypass_gate_3v256x8m81_7/m3_n41_5682# ypass_gate_3v256x8m81_7/m3_n41_6881#
Xypass_gate_3v256x8m81_1 ypass_gate_3v256x8m81_7/vss ypass_gate_3v256x8m81_7/vdd ypass_gate_3v256x8m81_1/b
+ ypass_gate_3v256x8m81_1/bb ypass_gate_3v256x8m81_1/ypass ypass_gate_3v256x8m81_7/pcb
+ ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_7/m3_n41_6881# ypass_gate_3v256x8m81_7/m3_n41_5924#
+ ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_1/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5682# ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5440#
+ ypass_gate_3v256x8m81_7/m3_n41_6156# VSUBS ypass_gate_3v256x8m81_1/db ypass_gate_3v256x8m81
Xypass_gate_3v256x8m81_2 ypass_gate_3v256x8m81_7/vss ypass_gate_3v256x8m81_7/vdd ypass_gate_3v256x8m81_2/b
+ ypass_gate_3v256x8m81_2/bb ypass_gate_3v256x8m81_2/ypass ypass_gate_3v256x8m81_7/pcb
+ ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_7/m3_n41_6881# ypass_gate_3v256x8m81_7/m3_n41_5924#
+ ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_2/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5682# ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5440#
+ ypass_gate_3v256x8m81_7/m3_n41_6156# VSUBS ypass_gate_3v256x8m81_4/db ypass_gate_3v256x8m81
Xypass_gate_3v256x8m81_3 ypass_gate_3v256x8m81_7/vss ypass_gate_3v256x8m81_7/vdd ypass_gate_3v256x8m81_3/b
+ ypass_gate_3v256x8m81_3/bb ypass_gate_3v256x8m81_3/ypass ypass_gate_3v256x8m81_7/pcb
+ ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_7/m3_n41_6881# ypass_gate_3v256x8m81_7/m3_n41_5924#
+ ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_3/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5682# ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5440#
+ ypass_gate_3v256x8m81_7/m3_n41_6156# VSUBS ypass_gate_3v256x8m81_5/db ypass_gate_3v256x8m81
Xypass_gate_3v256x8m81_4 ypass_gate_3v256x8m81_7/vss ypass_gate_3v256x8m81_7/vdd ypass_gate_3v256x8m81_4/b
+ ypass_gate_3v256x8m81_4/bb ypass_gate_3v256x8m81_4/ypass ypass_gate_3v256x8m81_7/pcb
+ ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_7/m3_n41_6881# ypass_gate_3v256x8m81_7/m3_n41_5924#
+ ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_4/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5682# ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5440#
+ ypass_gate_3v256x8m81_7/m3_n41_6156# VSUBS ypass_gate_3v256x8m81_4/db ypass_gate_3v256x8m81
Xypass_gate_3v256x8m81_5 ypass_gate_3v256x8m81_7/vss ypass_gate_3v256x8m81_7/vdd ypass_gate_3v256x8m81_5/b
+ ypass_gate_3v256x8m81_5/bb ypass_gate_3v256x8m81_5/ypass ypass_gate_3v256x8m81_7/pcb
+ ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_7/m3_n41_6881# ypass_gate_3v256x8m81_7/m3_n41_5924#
+ ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_5/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5682# ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5440#
+ ypass_gate_3v256x8m81_7/m3_n41_6156# VSUBS ypass_gate_3v256x8m81_5/db ypass_gate_3v256x8m81
Xypass_gate_3v256x8m81_6 ypass_gate_3v256x8m81_7/vss ypass_gate_3v256x8m81_7/vdd ypass_gate_3v256x8m81_6/b
+ ypass_gate_3v256x8m81_6/bb ypass_gate_3v256x8m81_6/ypass ypass_gate_3v256x8m81_7/pcb
+ ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_7/m3_n41_6881# ypass_gate_3v256x8m81_7/m3_n41_5924#
+ ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_6/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5682# ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5440#
+ ypass_gate_3v256x8m81_7/m3_n41_6156# VSUBS ypass_gate_3v256x8m81_7/db ypass_gate_3v256x8m81
Xypass_gate_3v256x8m81_7 ypass_gate_3v256x8m81_7/vss ypass_gate_3v256x8m81_7/vdd ypass_gate_3v256x8m81_7/b
+ ypass_gate_3v256x8m81_7/bb ypass_gate_3v256x8m81_7/ypass ypass_gate_3v256x8m81_7/pcb
+ ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_7/m3_n41_6881# ypass_gate_3v256x8m81_7/m3_n41_5924#
+ ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_7/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5682# ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5440#
+ ypass_gate_3v256x8m81_7/m3_n41_6156# VSUBS ypass_gate_3v256x8m81_7/db ypass_gate_3v256x8m81
Xypass_gate_a_3v256x8m81_0 ypass_gate_3v256x8m81_7/vss ypass_gate_a_3v256x8m81_0/b
+ ypass_gate_a_3v256x8m81_0/bb ypass_gate_a_3v256x8m81_0/ypass ypass_gate_3v256x8m81_7/pcb
+ ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_7/m3_n41_6881# ypass_gate_3v256x8m81_7/m3_n41_5924#
+ ypass_gate_3v256x8m81_7/m3_n41_6639# ypass_gate_3v256x8m81_7/vdd_uq0 ypass_gate_3v256x8m81_7/m3_n41_5682#
+ ypass_gate_3v256x8m81_7/vdd ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ VSUBS ypass_gate_3v256x8m81_1/db ypass_gate_a_3v256x8m81_0/pmos_1p2$$46889004_3v256x8m81_1/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_7/m3_n41_5198# ypass_gate_3v256x8m81_7/m3_n41_5440# ypass_gate_3v256x8m81_7/m3_n41_6156#
+ ypass_gate_a_3v256x8m81
.ends

.subckt pmos_5p04310591302018_3v256x8m81 D_uq1 a_20_n45# D_uq0 D a_181_n45# S_uq2
+ a_502_n45# S_uq1 a_662_n45# a_n140_n45# S_uq0 S a_341_n45# w_n314_n86#
X0 S a_341_n45# D w_n314_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
X1 S_uq0 a_662_n45# D_uq0 w_n314_n86# pfet_03v3 ad=0.4642p pd=2.99u as=0.2743p ps=1.575u w=1.055u l=0.28u
X2 D_uq0 a_502_n45# S w_n314_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.27692p ps=1.58u w=1.055u l=0.28u
X3 S_uq1 a_20_n45# D_uq1 w_n314_n86# pfet_03v3 ad=0.27692p pd=1.58u as=0.2743p ps=1.575u w=1.055u l=0.28u
X4 D a_181_n45# S_uq1 w_n314_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.27692p ps=1.58u w=1.055u l=0.28u
X5 D_uq1 a_n140_n45# S_uq2 w_n314_n86# pfet_03v3 ad=0.2743p pd=1.575u as=0.4642p ps=2.99u w=1.055u l=0.28u
.ends

.subckt pmos_1p2$$46549036_3v256x8m81 a_327_n34# w_n188_n50# pmos_5p04310591302018_3v256x8m81_0/D_uq1
+ pmos_5p04310591302018_3v256x8m81_0/D_uq0 pmos_5p04310591302018_3v256x8m81_0/S a_488_n34#
+ a_n154_n34# a_167_n34# pmos_5p04310591302018_3v256x8m81_0/D a_6_n34# pmos_5p04310591302018_3v256x8m81_0/S_uq2
+ pmos_5p04310591302018_3v256x8m81_0/S_uq1 a_648_n34# pmos_5p04310591302018_3v256x8m81_0/S_uq0
Xpmos_5p04310591302018_3v256x8m81_0 pmos_5p04310591302018_3v256x8m81_0/D_uq1 a_6_n34#
+ pmos_5p04310591302018_3v256x8m81_0/D_uq0 pmos_5p04310591302018_3v256x8m81_0/D a_167_n34#
+ pmos_5p04310591302018_3v256x8m81_0/S_uq2 a_488_n34# pmos_5p04310591302018_3v256x8m81_0/S_uq1
+ a_648_n34# a_n154_n34# pmos_5p04310591302018_3v256x8m81_0/S_uq0 pmos_5p04310591302018_3v256x8m81_0/S
+ a_327_n34# w_n188_n50# pmos_5p04310591302018_3v256x8m81
.ends

.subckt pmos_5p04310591302021_3v256x8m81 a_76_n44# D_uq0 D a_n84_n44# w_n258_n86#
+ S_uq1 S_uq0 S a_237_n44# a_397_n44#
X0 S_uq0 a_397_n44# D_uq0 w_n258_n86# pfet_03v3 ad=0.1848p pd=1.72u as=0.1092p ps=0.94u w=0.42u l=0.28u
X1 D_uq0 a_237_n44# S w_n258_n86# pfet_03v3 ad=0.1092p pd=0.94u as=0.11025p ps=0.945u w=0.42u l=0.28u
X2 D a_n84_n44# S_uq1 w_n258_n86# pfet_03v3 ad=0.1092p pd=0.94u as=0.1848p ps=1.72u w=0.42u l=0.28u
X3 S a_76_n44# D w_n258_n86# pfet_03v3 ad=0.11025p pd=0.945u as=0.1092p ps=0.94u w=0.42u l=0.28u
.ends

.subckt pmos_1p2$$46896172_3v256x8m81 w_n133_n66# pmos_5p04310591302021_3v256x8m81_0/D_uq0
+ pmos_5p04310591302021_3v256x8m81_0/S pmos_5p04310591302021_3v256x8m81_0/a_n84_n44#
+ pmos_5p04310591302021_3v256x8m81_0/D pmos_5p04310591302021_3v256x8m81_0/S_uq1 pmos_5p04310591302021_3v256x8m81_0/a_76_n44#
+ pmos_5p04310591302021_3v256x8m81_0/S_uq0 pmos_5p04310591302021_3v256x8m81_0/a_237_n44#
+ pmos_5p04310591302021_3v256x8m81_0/a_397_n44#
Xpmos_5p04310591302021_3v256x8m81_0 pmos_5p04310591302021_3v256x8m81_0/a_76_n44# pmos_5p04310591302021_3v256x8m81_0/D_uq0
+ pmos_5p04310591302021_3v256x8m81_0/D pmos_5p04310591302021_3v256x8m81_0/a_n84_n44#
+ w_n133_n66# pmos_5p04310591302021_3v256x8m81_0/S_uq1 pmos_5p04310591302021_3v256x8m81_0/S_uq0
+ pmos_5p04310591302021_3v256x8m81_0/S pmos_5p04310591302021_3v256x8m81_0/a_237_n44#
+ pmos_5p04310591302021_3v256x8m81_0/a_397_n44# pmos_5p04310591302021_3v256x8m81
.ends

.subckt pmos_1p2$$46897196_3v256x8m81 w_n133_n66# a_n42_n34# pmos_5p04310591302020_3v256x8m81_0/D
+ pmos_5p04310591302020_3v256x8m81_0/S_uq0 a_118_n34# pmos_5p04310591302020_3v256x8m81_0/S
Xpmos_5p04310591302020_3v256x8m81_0 pmos_5p04310591302020_3v256x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302020_3v256x8m81_0/S_uq0 pmos_5p04310591302020_3v256x8m81_0/S
+ pmos_5p04310591302020_3v256x8m81
.ends

.subckt nmos_5p04310591302015_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.6996p pd=4.06u as=0.6996p ps=4.06u w=1.59u l=0.28u
.ends

.subckt nmos_1p2$$46553132_3v256x8m81 nmos_5p04310591302015_3v256x8m81_0/S a_n14_n34#
+ nmos_5p04310591302015_3v256x8m81_0/D VSUBS
Xnmos_5p04310591302015_3v256x8m81_0 nmos_5p04310591302015_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302015_3v256x8m81_0/S VSUBS nmos_5p04310591302015_3v256x8m81
.ends

.subckt nmos_1p2$$45107244_3v256x8m81 nmos_5p04310591302012_3v256x8m81_0/S_uq1 a_223_n34#
+ nmos_5p04310591302012_3v256x8m81_0/S_uq0 a_383_n34# nmos_5p04310591302012_3v256x8m81_0/S
+ nmos_5p04310591302012_3v256x8m81_0/D_uq0 a_n96_n34# a_63_n34# nmos_5p04310591302012_3v256x8m81_0/D
+ VSUBS
Xnmos_5p04310591302012_3v256x8m81_0 a_n96_n34# nmos_5p04310591302012_3v256x8m81_0/D_uq0
+ nmos_5p04310591302012_3v256x8m81_0/D a_63_n34# nmos_5p04310591302012_3v256x8m81_0/S_uq1
+ nmos_5p04310591302012_3v256x8m81_0/S_uq0 nmos_5p04310591302012_3v256x8m81_0/S a_223_n34#
+ a_383_n34# VSUBS nmos_5p04310591302012_3v256x8m81
.ends

.subckt nmos_5p04310591302016_3v256x8m81 D_uq2 a_124_n45# D_uq1 a_284_n45# D_uq0 D
+ a_446_n45# a_768_n45# a_n198_n45# a_n38_n45# S_uq2 S_uq3 S_uq1 S_uq0 a_606_n45#
+ S a_928_n45# VSUBS
X0 S_uq0 a_928_n45# D_uq0 VSUBS nfet_03v3 ad=0.7155p pd=4.08u as=0.4134p ps=2.11u w=1.59u l=0.28u
X1 D_uq2 a_n198_n45# S_uq3 VSUBS nfet_03v3 ad=0.4134p pd=2.11u as=0.70755p ps=4.07u w=1.59u l=0.28u
X2 S_uq2 a_n38_n45# D_uq2 VSUBS nfet_03v3 ad=0.42135p pd=2.12u as=0.4134p ps=2.11u w=1.59u l=0.28u
X3 S a_606_n45# D VSUBS nfet_03v3 ad=0.42135p pd=2.12u as=0.4134p ps=2.11u w=1.59u l=0.28u
X4 D_uq0 a_768_n45# S VSUBS nfet_03v3 ad=0.4134p pd=2.11u as=0.42135p ps=2.12u w=1.59u l=0.28u
X5 D a_446_n45# S_uq1 VSUBS nfet_03v3 ad=0.4134p pd=2.11u as=0.42135p ps=2.12u w=1.59u l=0.28u
X6 S_uq1 a_284_n45# D_uq1 VSUBS nfet_03v3 ad=0.42135p pd=2.12u as=0.4134p ps=2.11u w=1.59u l=0.28u
X7 D_uq1 a_124_n45# S_uq2 VSUBS nfet_03v3 ad=0.4134p pd=2.11u as=0.42135p ps=2.12u w=1.59u l=0.28u
.ends

.subckt nmos_1p2$$46552108_3v256x8m81 nmos_5p04310591302016_3v256x8m81_0/D_uq2 nmos_5p04310591302016_3v256x8m81_0/D_uq1
+ nmos_5p04310591302016_3v256x8m81_0/D_uq0 nmos_5p04310591302016_3v256x8m81_0/a_124_n45#
+ nmos_5p04310591302016_3v256x8m81_0/a_284_n45# nmos_5p04310591302016_3v256x8m81_0/a_446_n45#
+ nmos_5p04310591302016_3v256x8m81_0/a_768_n45# nmos_5p04310591302016_3v256x8m81_0/a_n38_n45#
+ nmos_5p04310591302016_3v256x8m81_0/S nmos_5p04310591302016_3v256x8m81_0/S_uq3 nmos_5p04310591302016_3v256x8m81_0/S_uq2
+ nmos_5p04310591302016_3v256x8m81_0/a_n198_n45# nmos_5p04310591302016_3v256x8m81_0/S_uq1
+ nmos_5p04310591302016_3v256x8m81_0/S_uq0 nmos_5p04310591302016_3v256x8m81_0/a_606_n45#
+ nmos_5p04310591302016_3v256x8m81_0/a_928_n45# nmos_5p04310591302016_3v256x8m81_0/D
+ VSUBS
Xnmos_5p04310591302016_3v256x8m81_0 nmos_5p04310591302016_3v256x8m81_0/D_uq2 nmos_5p04310591302016_3v256x8m81_0/a_124_n45#
+ nmos_5p04310591302016_3v256x8m81_0/D_uq1 nmos_5p04310591302016_3v256x8m81_0/a_284_n45#
+ nmos_5p04310591302016_3v256x8m81_0/D_uq0 nmos_5p04310591302016_3v256x8m81_0/D nmos_5p04310591302016_3v256x8m81_0/a_446_n45#
+ nmos_5p04310591302016_3v256x8m81_0/a_768_n45# nmos_5p04310591302016_3v256x8m81_0/a_n198_n45#
+ nmos_5p04310591302016_3v256x8m81_0/a_n38_n45# nmos_5p04310591302016_3v256x8m81_0/S_uq2
+ nmos_5p04310591302016_3v256x8m81_0/S_uq3 nmos_5p04310591302016_3v256x8m81_0/S_uq1
+ nmos_5p04310591302016_3v256x8m81_0/S_uq0 nmos_5p04310591302016_3v256x8m81_0/a_606_n45#
+ nmos_5p04310591302016_3v256x8m81_0/S nmos_5p04310591302016_3v256x8m81_0/a_928_n45#
+ VSUBS nmos_5p04310591302016_3v256x8m81
.ends

.subckt pmos_5p04310591302019_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.1848p pd=1.72u as=0.1848p ps=1.72u w=0.42u l=0.28u
.ends

.subckt pmos_1p2$$46898220_3v256x8m81 w_n133_n66# a_n14_84# pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_5p04310591302019_3v256x8m81_0/D
Xpmos_5p04310591302019_3v256x8m81_0 pmos_5p04310591302019_3v256x8m81_0/D a_n14_84#
+ w_n133_n66# pmos_5p04310591302019_3v256x8m81_0/S pmos_5p04310591302019_3v256x8m81
.ends

.subckt nmos_5p04310591302017_3v256x8m81 D_uq2 D_uq1 a_n37_n44# D_uq0 D a_929_n44#
+ a_125_n44# a_285_n44# a_447_n44# a_769_n44# S_uq2 S_uq3 S_uq1 S_uq0 S a_607_n44#
+ a_n197_n44# VSUBS
X0 D_uq0 a_769_n44# S VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.35112p ps=1.855u w=1.325u l=0.28u
X1 D a_447_n44# S_uq1 VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.35112p ps=1.855u w=1.325u l=0.28u
X2 D_uq2 a_n197_n44# S_uq3 VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.583p ps=3.53u w=1.325u l=0.28u
X3 S_uq2 a_n37_n44# D_uq2 VSUBS nfet_03v3 ad=0.35112p pd=1.855u as=0.3445p ps=1.845u w=1.325u l=0.28u
X4 S_uq1 a_285_n44# D_uq1 VSUBS nfet_03v3 ad=0.35112p pd=1.855u as=0.3445p ps=1.845u w=1.325u l=0.28u
X5 D_uq1 a_125_n44# S_uq2 VSUBS nfet_03v3 ad=0.3445p pd=1.845u as=0.35112p ps=1.855u w=1.325u l=0.28u
X6 S_uq0 a_929_n44# D_uq0 VSUBS nfet_03v3 ad=0.58963p pd=3.54u as=0.3445p ps=1.845u w=1.325u l=0.28u
X7 S a_607_n44# D VSUBS nfet_03v3 ad=0.35112p pd=1.855u as=0.3445p ps=1.845u w=1.325u l=0.28u
.ends

.subckt nmos_1p2$$46550060_3v256x8m81 nmos_5p04310591302017_3v256x8m81_0/D_uq2 nmos_5p04310591302017_3v256x8m81_0/D_uq1
+ nmos_5p04310591302017_3v256x8m81_0/D nmos_5p04310591302017_3v256x8m81_0/D_uq0 a_915_n34#
+ a_111_n34# a_271_n34# a_433_n34# a_593_n34# a_n51_n34# a_755_n34# nmos_5p04310591302017_3v256x8m81_0/S_uq3
+ a_n210_n34# nmos_5p04310591302017_3v256x8m81_0/S_uq1 nmos_5p04310591302017_3v256x8m81_0/S_uq2
+ nmos_5p04310591302017_3v256x8m81_0/S nmos_5p04310591302017_3v256x8m81_0/S_uq0 VSUBS
Xnmos_5p04310591302017_3v256x8m81_0 nmos_5p04310591302017_3v256x8m81_0/D_uq2 nmos_5p04310591302017_3v256x8m81_0/D_uq1
+ a_n51_n34# nmos_5p04310591302017_3v256x8m81_0/D_uq0 nmos_5p04310591302017_3v256x8m81_0/D
+ a_915_n34# a_111_n34# a_271_n34# a_433_n34# a_755_n34# nmos_5p04310591302017_3v256x8m81_0/S_uq2
+ nmos_5p04310591302017_3v256x8m81_0/S_uq3 nmos_5p04310591302017_3v256x8m81_0/S_uq1
+ nmos_5p04310591302017_3v256x8m81_0/S_uq0 nmos_5p04310591302017_3v256x8m81_0/S a_593_n34#
+ a_n210_n34# VSUBS nmos_5p04310591302017_3v256x8m81
.ends

.subckt nmos_1p2$$46551084_3v256x8m81 nmos_5p04310591302010_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v256x8m81_0/S VSUBS
Xnmos_5p04310591302010_3v256x8m81_0 nmos_5p04310591302010_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v256x8m81_0/S VSUBS nmos_5p04310591302010_3v256x8m81
.ends

.subckt sa_3v256x8m81 qp qn wep se pcb db pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D
+ vdd d vss
Xpmos_1p2$$46549036_3v256x8m81_0 nmos_1p2$$46551084_3v256x8m81_0/nmos_5p04310591302010_3v256x8m81_0/S
+ vdd qn nmos_1p2$$46551084_3v256x8m81_0/nmos_5p04310591302010_3v256x8m81_0/S vdd
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D
+ nmos_1p2$$46551084_3v256x8m81_0/nmos_5p04310591302010_3v256x8m81_0/S qp pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D
+ vdd vdd pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S vdd
+ pmos_1p2$$46549036_3v256x8m81
Xpmos_1p2$$46896172_3v256x8m81_0 pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D
+ pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D pmos_1p2$$46896172_3v256x8m81
Xpmos_1p2$$46897196_3v256x8m81_0 pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D
+ se pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S d se d pmos_1p2$$46897196_3v256x8m81
Xpmos_1p2$$46897196_3v256x8m81_1 pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D
+ se pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D db se db
+ pmos_1p2$$46897196_3v256x8m81
Xpmos_1p2$$46897196_3v256x8m81_2 pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D
+ se pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D db se db
+ pmos_1p2$$46897196_3v256x8m81
Xpmos_1p2$$46897196_3v256x8m81_3 pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D
+ se pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S d se d pmos_1p2$$46897196_3v256x8m81
Xnmos_1p2$$46553132_3v256x8m81_0 pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D
+ vss vss vss nmos_1p2$$46553132_3v256x8m81
Xnmos_1p2$$46553132_3v256x8m81_1 vss vss pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D
+ vss nmos_1p2$$46553132_3v256x8m81
Xnmos_1p2$$45107244_3v256x8m81_0 qn nmos_1p2$$46551084_3v256x8m81_0/nmos_5p04310591302010_3v256x8m81_0/S
+ qp nmos_1p2$$46551084_3v256x8m81_0/nmos_5p04310591302010_3v256x8m81_0/S qp vss pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D
+ nmos_1p2$$46551084_3v256x8m81_0/nmos_5p04310591302010_3v256x8m81_0/S vss vss nmos_1p2$$45107244_3v256x8m81
Xnmos_1p2$$46552108_3v256x8m81_0 nmos_1p2$$46552108_3v256x8m81_0/nmos_5p04310591302016_3v256x8m81_0/D
+ nmos_1p2$$46552108_3v256x8m81_0/nmos_5p04310591302016_3v256x8m81_0/D nmos_1p2$$46552108_3v256x8m81_0/nmos_5p04310591302016_3v256x8m81_0/D
+ pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D
+ pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D
+ pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S nmos_1p2$$46552108_3v256x8m81_0/nmos_5p04310591302016_3v256x8m81_0/D
+ vss nmos_1p2$$46552108_3v256x8m81
Xpmos_1p2$$46898220_3v256x8m81_0 pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S pmos_1p2$$46898220_3v256x8m81
Xpmos_1p2$$46898220_3v256x8m81_1 pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D pmos_1p2$$46898220_3v256x8m81
Xnmos_1p2$$46550060_3v256x8m81_0 nmos_1p2$$46552108_3v256x8m81_0/nmos_5p04310591302016_3v256x8m81_0/D
+ nmos_1p2$$46552108_3v256x8m81_0/nmos_5p04310591302016_3v256x8m81_0/D nmos_1p2$$46552108_3v256x8m81_0/nmos_5p04310591302016_3v256x8m81_0/D
+ nmos_1p2$$46552108_3v256x8m81_0/nmos_5p04310591302016_3v256x8m81_0/D se se se se
+ se se se vss se vss vss vss vss vss nmos_1p2$$46550060_3v256x8m81
Xpmos_1p2$$46286892_3v256x8m81_0 pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D
+ db d pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D pcb pcb
+ pcb pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D pmos_1p2$$46286892_3v256x8m81
Xpmos_1p2$$46285868_3v256x8m81_0 pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/D
+ pmos_1p2$$46897196_3v256x8m81_2/pmos_5p04310591302020_3v256x8m81_0/D pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ pcb pmos_1p2$$46285868_3v256x8m81
Xnmos_1p2$$46551084_3v256x8m81_0 vss pmos_1p2$$46898220_3v256x8m81_1/pmos_5p04310591302019_3v256x8m81_0/S
+ nmos_1p2$$46551084_3v256x8m81_0/nmos_5p04310591302010_3v256x8m81_0/S vss nmos_1p2$$46551084_3v256x8m81
.ends

.subckt saout_R_m2_3v256x8m81 ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] GWEN datain
+ b[5] b[4] b[2] b[1] b[0] bb[6] q bb[3] bb[0] bb[1] pcb vss_uq6 vdd_uq0 vdd_uq2 vdd_uq4
+ vdd_uq6 pcb_uq0 datain_uq0 mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ bb[5] sa_3v256x8m81_0/pcb sa_3v256x8m81_0/d mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ GWE bb[2] WEN mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb b[3] ypass[7] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass b[6] bb[4] vdd mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ din_3v256x8m81_0/men mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass bb[7] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ vdd_uq3 ypass[1] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass b[7] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass
+ vss mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass vdd_uq1 vdd_uq5 sacntl_2_3v256x8m81_0/vdd_uq0
Xsacntl_2_3v256x8m81_0 sa_3v256x8m81_0/pcb sa_3v256x8m81_0/se sacntl_2_3v256x8m81_0/vdd_uq0
+ sacntl_2_3v256x8m81_0/pmos_5p04310591302027_3v256x8m81_1/S_uq0 sacntl_2_3v256x8m81_0/pmos_5p04310591302027_3v256x8m81_2/S_uq0
+ din_3v256x8m81_0/men vdd_uq0 vss sacntl_2_3v256x8m81
Xoutbuf_oe_3v256x8m81_0 sa_3v256x8m81_0/qp sa_3v256x8m81_0/qn sa_3v256x8m81_0/se q
+ GWE vdd_uq3 vss outbuf_oe_3v256x8m81
Xdin_3v256x8m81_0 vss datain din_3v256x8m81_0/men sa_3v256x8m81_0/db sa_3v256x8m81_0/d
+ sa_3v256x8m81_0/wep vdd_uq5 vdd_uq3 sa_3v256x8m81_0/pcb vss din_3v256x8m81
Xwen_wm1_3v256x8m81_0 GWEN din_3v256x8m81_0/men sa_3v256x8m81_0/wep vss vdd WEN vdd_uq1
+ wen_wm1_3v256x8m81
Xmux821_3v256x8m81_0 sa_3v256x8m81_0/d mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ bb[5] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb b[6] mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ sa_3v256x8m81_0/db mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass sa_3v256x8m81_0/d
+ sa_3v256x8m81_0/d mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/ypass ypass[7] b[3] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ bb[2] sa_3v256x8m81_0/db sa_3v256x8m81_0/db sa_3v256x8m81_0/d sa_3v256x8m81_0/d
+ bb[7] sa_3v256x8m81_0/d mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass
+ sa_3v256x8m81_0/pcb ypass[7] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ b[7] ypass[1] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ bb[4] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b sa_3v256x8m81_0/d mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass
+ sa_3v256x8m81_0/d vss sa_3v256x8m81_0/db mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/ypass
+ mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass mux821_3v256x8m81
Xsa_3v256x8m81_0 sa_3v256x8m81_0/qp sa_3v256x8m81_0/qn sa_3v256x8m81_0/wep sa_3v256x8m81_0/se
+ sa_3v256x8m81_0/pcb sa_3v256x8m81_0/db vdd_uq5 vdd_uq3 sa_3v256x8m81_0/d vss sa_3v256x8m81
.ends

.subckt x018SRAM_cell1_2x_3v256x8m81 018SRAM_cell1_3v256x8m81_0/m3_82_330# 018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# 018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_3v256x8m81_0/a_62_178# 018SRAM_cell1_3v256x8m81_0/w_30_512# 018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_3v256x8m81_1/a_62_178# VSUBS
X018SRAM_cell1_3v256x8m81_0 018SRAM_cell1_3v256x8m81_0/m3_82_330# 018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_3v256x8m81_0/a_62_178# 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_3v256x8m81_1/a_110_96# VSUBS
+ x018SRAM_cell1_3v256x8m81
X018SRAM_cell1_3v256x8m81_1 018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_3v256x8m81_1/a_62_178# 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_3v256x8m81_1/a_110_96# VSUBS
+ x018SRAM_cell1_3v256x8m81
.ends

.subckt Cell_array8x8_3v256x8m81 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96# VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
X018SRAM_cell1_2x_3v256x8m81_0[0|0] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[1|0] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[2|0] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[3|0] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[4|0] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[5|0] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[6|0] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[7|0] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[8|0] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[9|0] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[10|0] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[11|0] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[12|0] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[13|0] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[14|0] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[15|0] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[0|1] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[1|1] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[2|1] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[3|1] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[4|1] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[5|1] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[6|1] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[7|1] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[8|1] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[9|1] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[10|1] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[11|1] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[12|1] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[13|1] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[14|1] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[15|1] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[0|2] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[1|2] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[2|2] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[3|2] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[4|2] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[5|2] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[6|2] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[7|2] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[8|2] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[9|2] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[10|2] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[11|2] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[12|2] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[13|2] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[14|2] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[15|2] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[0|3] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[1|3] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[2|3] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[3|3] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[4|3] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[5|3] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[6|3] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[7|3] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[8|3] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[9|3] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[10|3] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[11|3] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[12|3] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[13|3] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[14|3] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[15|3] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[0|4] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[1|4] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[2|4] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[3|4] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[4|4] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[5|4] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[6|4] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[7|4] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[8|4] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[9|4] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[10|4] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[11|4] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[12|4] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[13|4] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[14|4] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[15|4] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[0|5] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[1|5] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[2|5] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[3|5] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[4|5] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[5|5] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[6|5] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[7|5] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[8|5] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[9|5] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[10|5] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[11|5] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[12|5] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[13|5] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[14|5] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[15|5] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[0|6] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[1|6] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[2|6] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[3|6] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[4|6] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[5|6] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[6|6] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[7|6] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[8|6] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[9|6] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[10|6] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[11|6] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[12|6] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[13|6] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[14|6] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[15|6] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[0|7] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[1|7] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[2|7] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[3|7] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[4|7] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[5|7] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[6|7] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[7|7] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[8|7] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[9|7] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[10|7] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[11|7] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[12|7] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[13|7] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[14|7] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0[15|7] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_0[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[0|0] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[1|0] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[2|0] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[3|0] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[4|0] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[5|0] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[6|0] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[7|0] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[8|0] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[9|0] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[10|0] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[11|0] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[12|0] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[13|0] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[14|0] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[15|0] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[0|1] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[1|1] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[2|1] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[3|1] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[4|1] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[5|1] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[6|1] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[7|1] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[8|1] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[9|1] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[10|1] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[11|1] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[12|1] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[13|1] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[14|1] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[15|1] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[0|2] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[1|2] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[2|2] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[3|2] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[4|2] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[5|2] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[6|2] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[7|2] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[8|2] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[9|2] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[10|2] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[11|2] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[12|2] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[13|2] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[14|2] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[15|2] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[0|3] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[1|3] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[2|3] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[3|3] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[4|3] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[5|3] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[6|3] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[7|3] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[8|3] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[9|3] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[10|3] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[11|3] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[12|3] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[13|3] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[14|3] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[15|3] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[0|4] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[1|4] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[2|4] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[3|4] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[4|4] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[5|4] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[6|4] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[7|4] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[8|4] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[9|4] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[10|4] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[11|4] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[12|4] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[13|4] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[14|4] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[15|4] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[0|5] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[1|5] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[2|5] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[3|5] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[4|5] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[5|5] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[6|5] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[7|5] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[8|5] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[9|5] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[10|5] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[11|5] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[12|5] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[13|5] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[14|5] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[15|5] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[0|6] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[1|6] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[2|6] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[3|6] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[4|6] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[5|6] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[6|6] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[7|6] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[8|6] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[9|6] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[10|6] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[11|6] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[12|6] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[13|6] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[14|6] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[15|6] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[0|7] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[1|7] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[2|7] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[3|7] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[4|7] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[5|7] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[6|7] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[7|7] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[8|7] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[9|7] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[10|7] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[11|7] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[12|7] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[13|7] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[14|7] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1[15|7] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_1[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[0|0] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[1|0] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[2|0] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[3|0] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[4|0] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[5|0] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[6|0] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[7|0] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[8|0] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[9|0] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[10|0] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[11|0] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[12|0] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[13|0] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[14|0] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[15|0] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[0|1] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[1|1] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[2|1] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[3|1] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[4|1] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[5|1] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[6|1] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[7|1] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[8|1] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[9|1] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[10|1] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[11|1] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[12|1] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[13|1] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[14|1] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[15|1] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[0|2] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[1|2] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[2|2] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[3|2] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[4|2] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[5|2] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[6|2] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[7|2] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[8|2] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[9|2] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[10|2] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[11|2] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[12|2] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[13|2] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[14|2] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[15|2] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[0|3] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[1|3] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[2|3] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[3|3] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[4|3] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[5|3] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[6|3] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[7|3] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[8|3] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[9|3] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[10|3] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[11|3] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[12|3] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[13|3] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[14|3] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[15|3] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[0|4] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[1|4] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[2|4] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[3|4] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[4|4] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[5|4] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[6|4] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[7|4] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[8|4] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[9|4] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[10|4] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[11|4] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[12|4] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[13|4] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[14|4] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[15|4] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[0|5] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[1|5] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[2|5] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[3|5] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[4|5] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[5|5] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[6|5] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[7|5] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[8|5] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[9|5] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[10|5] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[11|5] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[12|5] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[13|5] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[14|5] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[15|5] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[0|6] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[1|6] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[2|6] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[3|6] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[4|6] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[5|6] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[6|6] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[7|6] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[8|6] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[9|6] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[10|6] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[11|6] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[12|6] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[13|6] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[14|6] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[15|6] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[0|7] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[1|7] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[2|7] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[3|7] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[4|7] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[5|7] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[6|7] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[7|7] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[8|7] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[9|7] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[10|7] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[11|7] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[12|7] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[13|7] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[14|7] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2[15|7] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_2[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[0|0] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[1|0] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[2|0] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[3|0] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[4|0] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[5|0] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[6|0] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[7|0] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[8|0] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[9|0] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[10|0] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[11|0] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[12|0] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[13|0] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[14|0] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[15|0] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|0]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[0|1] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[1|1] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[2|1] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[3|1] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[4|1] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[5|1] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[6|1] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[7|1] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[8|1] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[9|1] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[10|1] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[11|1] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[12|1] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[13|1] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[14|1] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[15|1] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|1]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[0|2] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[1|2] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[2|2] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[3|2] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[4|2] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[5|2] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[6|2] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[7|2] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[8|2] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[9|2] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[10|2] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[11|2] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[12|2] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[13|2] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[14|2] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[15|2] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|2]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[0|3] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[1|3] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[2|3] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[3|3] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[4|3] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[5|3] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[6|3] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[7|3] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[8|3] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[9|3] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[10|3] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[11|3] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[12|3] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[13|3] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[14|3] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[15|3] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|3]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[0|4] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[1|4] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[2|4] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[3|4] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[4|4] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[5|4] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[6|4] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[7|4] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[8|4] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[9|4] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[10|4] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[11|4] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[12|4] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[13|4] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[14|4] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[15|4] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|4]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[0|5] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[1|5] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[2|5] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[3|5] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[4|5] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[5|5] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[6|5] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[7|5] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[8|5] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[9|5] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[10|5] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[11|5] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[12|5] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[13|5] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[14|5] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[15|5] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|5]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[0|6] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[1|6] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[2|6] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[3|6] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[4|6] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[5|6] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[6|6] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[7|6] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[8|6] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[9|6] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[10|6] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[11|6] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[12|6] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[13|6] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[14|6] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[15|6] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|6]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[0|7] 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[0]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[1|7] 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[1]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[2|7] 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[2]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[3|7] 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[3]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[4|7] 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[4]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[5|7] 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[5]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[6|7] 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[6]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[7|7] 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[7]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[8|7] 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[8]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[9|7] 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[10|7] 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[10]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[11|7] 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[11]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[12|7] 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[12]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[13|7] 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[13]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[14|7] 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[14]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3[15|7] 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ VSUBS 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_0/a_91_178#
+ 018SRAM_strap1_2x_3v256x8m81_3[9]/018SRAM_strap1_3v256x8m81_1/w_91_512# 018SRAM_cell1_2x_3v256x8m81_3[9|7]/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_strap1_2x_3v256x8m81_3[15]/018SRAM_strap1_3v256x8m81_1/a_91_178# VSUBS x018SRAM_cell1_2x_3v256x8m81
.ends

.subckt saout_m2_3v256x8m81 ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] GWEN GWE
+ bb[1] bb[4] bb[7] bb[6] b[5] b[7] b[2] datain q pcb vss_uq4 vdd vdd_uq0 vdd_uq1
+ vdd_uq2 pcb_uq0 pcb_uq1 b[2]_uq0 b[7]_uq0 b[5]_uq0 bb[6]_uq0 bb[7]_uq0 bb[5] bb[4]_uq0
+ bb[1]_uq0 mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ b[6] bb[2] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass WEN mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ b[4] din_3v256x8m81_0/men outbuf_oe_3v256x8m81_0/GWE mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ b[1] bb[3] ypass[7] vdd_uq4 mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass b[3]
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb VDD_uq0 mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass
+ vss mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ VDD vdd_uq3 VDD_uq1
Xsacntl_2_3v256x8m81_0 pcb_uq0 sa_3v256x8m81_0/se VDD_uq0 sacntl_2_3v256x8m81_0/pmos_5p04310591302027_3v256x8m81_1/S_uq0
+ sacntl_2_3v256x8m81_0/pmos_5p04310591302027_3v256x8m81_2/S_uq0 din_3v256x8m81_0/men
+ vdd_uq2 vss sacntl_2_3v256x8m81
Xoutbuf_oe_3v256x8m81_0 sa_3v256x8m81_0/qp sa_3v256x8m81_0/qn sa_3v256x8m81_0/se q
+ outbuf_oe_3v256x8m81_0/GWE vdd vss outbuf_oe_3v256x8m81
Xdin_3v256x8m81_0 vss datain din_3v256x8m81_0/men sa_3v256x8m81_0/db sa_3v256x8m81_0/d
+ sa_3v256x8m81_0/wep vdd_uq3 vdd pcb_uq0 vss din_3v256x8m81
Xwen_wm1_3v256x8m81_0 GWEN din_3v256x8m81_0/men sa_3v256x8m81_0/wep vss VDD_uq1 WEN
+ VDD wen_wm1_3v256x8m81
Xmux821_3v256x8m81_0 sa_3v256x8m81_0/d b[6] mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb bb[2] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ b[1] mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ sa_3v256x8m81_0/db mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass sa_3v256x8m81_0/d
+ sa_3v256x8m81_0/d mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass
+ ypass[7] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass b[4] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ bb[5] sa_3v256x8m81_0/db sa_3v256x8m81_0/db sa_3v256x8m81_0/d sa_3v256x8m81_0/d
+ mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb sa_3v256x8m81_0/d mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass pcb_uq0 ypass[7] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass
+ b[3] vdd_uq4 vdd_uq0 mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ bb[3] mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b sa_3v256x8m81_0/d mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ sa_3v256x8m81_0/d vss sa_3v256x8m81_0/db mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass
+ mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass mux821_3v256x8m81
Xsa_3v256x8m81_0 sa_3v256x8m81_0/qp sa_3v256x8m81_0/qn sa_3v256x8m81_0/wep sa_3v256x8m81_0/se
+ pcb_uq0 sa_3v256x8m81_0/db vdd_uq3 vdd sa_3v256x8m81_0/d vss sa_3v256x8m81
.ends

.subckt col_256a_3v256x8m81 ypass[0] ypass[1] ypass[3] ypass[4] ypass[5] ypass[7]
+ VDD WL[32] WL[31] WL[30] WL[20] WL[11] WL[10] WL[7] WL[18] WL[17] WL[16] WL[15]
+ WL[14] WL[13] WL[27] WL[26] ypass[6] ypass[2] b[1] b[7] b[10] b[13] b[16] b[22]
+ b[28] din[1] din[3] din[2] din[0] q[0] q[1] q[2] q[3] b[29] b[23] b[20] b[14] b[11]
+ b[8] bb[0] bb[1] bb[2] bb[8] bb[9] bb[11] bb[12] bb[13] bb[14] bb[15] bb[19] bb[21]
+ bb[22] bb[24] bb[26] bb[28] bb[29] bb[30] bb[31] b[30] b[27] b[0] b[3] b[18] pcb[0]
+ pcb[1] pcb[3] pcb[2] WEN[3] WEN[2] WEN[1] WEN[0] VDD_uq5 saout_R_m2_3v256x8m81_0/q
+ saout_R_m2_3v256x8m81_1/datain saout_m2_3v256x8m81_4/GWEN saout_m2_3v256x8m81_4/outbuf_oe_3v256x8m81_0/GWE
+ WL[1] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb saout_m2_3v256x8m81_4/q
+ WL[4] men saout_R_m2_3v256x8m81_0/vdd_uq4 saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ WL[21] m3_n771_22409# saout_R_m2_3v256x8m81_0/datain b[9] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ WL[24] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb saout_R_m2_3v256x8m81_0/GWE
+ VDD_uq4 saout_m2_3v256x8m81_3/b[6] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b b[25] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb WL[5] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ VDD_uq1 saout_m2_3v256x8m81_4/GWE saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ WL[8] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb saout_m2_3v256x8m81_3/b[1]
+ saout_R_m2_3v256x8m81_1/bb[5] WL[25] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_m2_3v256x8m81_4/b[6] saout_m2_3v256x8m81_3/bb[5] WL[2] WL[28] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ saout_R_m2_3v256x8m81_0/b[3] saout_m2_3v256x8m81_3/bb[3] saout_R_m2_3v256x8m81_1/q
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_3/q WL[22] saout_m2_3v256x8m81_4/b[3] saout_m2_3v256x8m81_4/datain
+ saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb b[31] saout_R_m2_3v256x8m81_1/GWE
+ saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b VDD_uq3 saout_m2_3v256x8m81_3/bb[2]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb VDD_uq2 WL[9]
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb bb[4] WL[12]
+ b[12] saout_m2_3v256x8m81_4/bb[5] GWE saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ WL[3] saout_m2_3v256x8m81_3/b[4] WL[29] b[5] WL[6] saout_R_m2_3v256x8m81_0/bb[4]
+ saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b saout_m2_3v256x8m81_3/datain
+ saout_R_m2_3v256x8m81_1/b[3] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ bb[17] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_1/b[6] saout_R_m2_3v256x8m81_1/bb[4] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_R_m2_3v256x8m81_0/bb[2] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ saout_m2_3v256x8m81_3/b[3] VDD_uq0 WL[23] saout_R_m2_3v256x8m81_1/bb[7] bb[10] VSS
+ WL[19] b[6] WL[0] bb[6]
Xsaout_R_m2_3v256x8m81_0 saout_R_m2_3v256x8m81_0/ypass[2] saout_R_m2_3v256x8m81_0/ypass[3]
+ saout_R_m2_3v256x8m81_0/ypass[4] saout_R_m2_3v256x8m81_0/ypass[5] saout_R_m2_3v256x8m81_0/ypass[6]
+ saout_m2_3v256x8m81_4/GWEN saout_R_m2_3v256x8m81_0/datain saout_R_m2_3v256x8m81_0/b[5]
+ saout_R_m2_3v256x8m81_0/b[4] saout_R_m2_3v256x8m81_0/b[2] saout_R_m2_3v256x8m81_0/b[1]
+ saout_R_m2_3v256x8m81_0/b[0] saout_R_m2_3v256x8m81_0/bb[6] saout_R_m2_3v256x8m81_0/q
+ saout_R_m2_3v256x8m81_0/bb[3] saout_R_m2_3v256x8m81_0/bb[0] saout_R_m2_3v256x8m81_0/bb[1]
+ saout_R_m2_3v256x8m81_0/pcb saout_R_m2_3v256x8m81_0/vss_uq6 VDD_uq2 saout_R_m2_3v256x8m81_0/vdd_uq2
+ saout_R_m2_3v256x8m81_0/vdd_uq4 saout_R_m2_3v256x8m81_0/vdd_uq6 saout_R_m2_3v256x8m81_0/pcb_uq0
+ saout_R_m2_3v256x8m81_0/datain_uq0 saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ bb[4] saout_R_m2_3v256x8m81_0/sa_3v256x8m81_0/pcb saout_R_m2_3v256x8m81_0/sa_3v256x8m81_0/d
+ saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b saout_R_m2_3v256x8m81_0/GWE
+ saout_R_m2_3v256x8m81_0/bb[2] WEN[0] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ saout_R_m2_3v256x8m81_0/b[3] ypass[5] ypass[2] ypass[0] b[5] saout_R_m2_3v256x8m81_0/bb[4]
+ VDD ypass[1] men saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b ypass[4] bb[6]
+ saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb VDD_uq3 VDD_uq5
+ ypass[6] b[6] ypass[3] VSS ypass[7] VDD_uq0 VDD_uq4 VDD_uq1 saout_R_m2_3v256x8m81
Xsaout_R_m2_3v256x8m81_1 saout_R_m2_3v256x8m81_1/ypass[2] saout_R_m2_3v256x8m81_1/ypass[3]
+ saout_R_m2_3v256x8m81_1/ypass[4] saout_R_m2_3v256x8m81_1/ypass[5] saout_R_m2_3v256x8m81_1/ypass[6]
+ saout_m2_3v256x8m81_4/GWEN saout_R_m2_3v256x8m81_1/datain saout_R_m2_3v256x8m81_1/b[5]
+ saout_R_m2_3v256x8m81_1/b[4] saout_R_m2_3v256x8m81_1/b[2] saout_R_m2_3v256x8m81_1/b[1]
+ saout_R_m2_3v256x8m81_1/b[0] saout_R_m2_3v256x8m81_1/bb[6] saout_R_m2_3v256x8m81_1/q
+ saout_R_m2_3v256x8m81_1/bb[3] saout_R_m2_3v256x8m81_1/bb[0] saout_R_m2_3v256x8m81_1/bb[1]
+ saout_R_m2_3v256x8m81_1/pcb saout_R_m2_3v256x8m81_1/vss_uq6 VDD_uq2 saout_R_m2_3v256x8m81_1/vdd_uq2
+ saout_R_m2_3v256x8m81_1/vdd_uq4 saout_R_m2_3v256x8m81_1/vdd_uq6 saout_R_m2_3v256x8m81_1/pcb_uq0
+ saout_R_m2_3v256x8m81_1/datain_uq0 saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_1/bb[5] saout_R_m2_3v256x8m81_1/sa_3v256x8m81_0/pcb saout_R_m2_3v256x8m81_1/sa_3v256x8m81_0/d
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b saout_R_m2_3v256x8m81_1/GWE
+ b[18] WEN[2] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ saout_R_m2_3v256x8m81_1/b[3] ypass[5] ypass[2] ypass[0] saout_R_m2_3v256x8m81_1/b[6]
+ saout_R_m2_3v256x8m81_1/bb[4] VDD ypass[1] men bb[17] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ ypass[4] saout_R_m2_3v256x8m81_1/bb[7] b[16] VDD_uq3 VDD_uq5 ypass[6] b[6] ypass[3]
+ VSS ypass[7] VDD_uq0 VDD_uq4 VDD_uq1 saout_R_m2_3v256x8m81
XCell_array8x8_3v256x8m81_0 saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b bb[8] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ b[10] saout_R_m2_3v256x8m81_0/b[3] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ bb[6] b[9] b[29] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb WL[22] bb[11]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb saout_R_m2_3v256x8m81_0/bb[4]
+ b[25] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b saout_R_m2_3v256x8m81_1/bb[4]
+ bb[10] bb[30] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ saout_m2_3v256x8m81_3/b[1] WL[28] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ WL[23] b[12] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ saout_m2_3v256x8m81_3/bb[3] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ WL[29] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b b[18] saout_m2_3v256x8m81_4/b[3]
+ b[31] b[16] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ saout_m2_3v256x8m81_3/bb[2] saout_m2_3v256x8m81_3/bb[5] saout_R_m2_3v256x8m81_1/b[6]
+ WL[24] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb saout_m2_3v256x8m81_4/bb[5]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_3/b[4] WL[10] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ WL[8] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb WL[17]
+ saout_R_m2_3v256x8m81_1/b[3] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ WL[0] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ WL[19] bb[17] bb[4] WL[9] WL[3] WL[6] saout_R_m2_3v256x8m81_0/bb[2] saout_m2_3v256x8m81_3/b[3]
+ WL[16] saout_m2_3v256x8m81_3/b[6] WL[1] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ WL[11] WL[21] saout_R_m2_3v256x8m81_1/bb[7] WL[31] WL[2] bb[24] saout_R_m2_3v256x8m81_1/bb[5]
+ WL[20] WL[12] WL[7] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ WL[5] WL[27] WL[25] WL[26] b[5] WL[30] WL[18] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ WL[15] WL[13] WL[4] saout_m2_3v256x8m81_4/b[6] VSS b[6] saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ WL[14] Cell_array8x8_3v256x8m81
Xsaout_m2_3v256x8m81_3 saout_m2_3v256x8m81_3/ypass[2] saout_m2_3v256x8m81_3/ypass[3]
+ saout_m2_3v256x8m81_3/ypass[4] saout_m2_3v256x8m81_3/ypass[5] saout_m2_3v256x8m81_3/ypass[6]
+ saout_m2_3v256x8m81_4/GWEN GWE saout_m2_3v256x8m81_3/bb[1] saout_m2_3v256x8m81_3/bb[4]
+ saout_m2_3v256x8m81_3/bb[7] saout_m2_3v256x8m81_3/bb[6] saout_m2_3v256x8m81_3/b[5]
+ saout_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/b[2] saout_m2_3v256x8m81_3/datain
+ saout_m2_3v256x8m81_3/q saout_m2_3v256x8m81_3/pcb saout_m2_3v256x8m81_3/vss_uq4
+ VDD_uq3 VDD_uq5 saout_m2_3v256x8m81_3/vdd_uq1 VDD_uq2 saout_m2_3v256x8m81_3/pcb_uq0
+ saout_m2_3v256x8m81_3/pcb_uq1 saout_m2_3v256x8m81_3/b[2]_uq0 saout_m2_3v256x8m81_3/b[7]_uq0
+ saout_m2_3v256x8m81_3/b[5]_uq0 saout_m2_3v256x8m81_3/bb[6]_uq0 saout_m2_3v256x8m81_3/bb[7]_uq0
+ saout_m2_3v256x8m81_3/bb[5] saout_m2_3v256x8m81_3/bb[4]_uq0 saout_m2_3v256x8m81_3/bb[1]_uq0
+ b[29] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_3/b[6] saout_m2_3v256x8m81_3/bb[2] ypass[2] WEN[3] b[31] bb[24]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb saout_m2_3v256x8m81_3/b[4]
+ men GWE b[25] ypass[0] bb[30] saout_m2_3v256x8m81_3/b[1] saout_m2_3v256x8m81_3/bb[3]
+ ypass[5] b[6] ypass[1] saout_m2_3v256x8m81_3/b[3] ypass[4] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb VDD_uq1 ypass[3]
+ VSS ypass[7] ypass[6] VDD_uq0 VDD_uq4 VDD saout_m2_3v256x8m81
Xsaout_m2_3v256x8m81_4 saout_m2_3v256x8m81_4/ypass[2] saout_m2_3v256x8m81_4/ypass[3]
+ saout_m2_3v256x8m81_4/ypass[4] saout_m2_3v256x8m81_4/ypass[5] saout_m2_3v256x8m81_4/ypass[6]
+ saout_m2_3v256x8m81_4/GWEN saout_m2_3v256x8m81_4/GWE saout_m2_3v256x8m81_4/bb[1]
+ saout_m2_3v256x8m81_4/bb[4] saout_m2_3v256x8m81_4/bb[7] saout_m2_3v256x8m81_4/bb[6]
+ saout_m2_3v256x8m81_4/b[5] saout_m2_3v256x8m81_4/b[7] saout_m2_3v256x8m81_4/b[2]
+ saout_m2_3v256x8m81_4/datain saout_m2_3v256x8m81_4/q saout_m2_3v256x8m81_4/pcb saout_m2_3v256x8m81_4/vss_uq4
+ VDD_uq3 VDD_uq5 saout_m2_3v256x8m81_4/vdd_uq1 VDD_uq2 saout_m2_3v256x8m81_4/pcb_uq0
+ saout_m2_3v256x8m81_4/pcb_uq1 saout_m2_3v256x8m81_4/b[2]_uq0 saout_m2_3v256x8m81_4/b[7]_uq0
+ saout_m2_3v256x8m81_4/b[5]_uq0 saout_m2_3v256x8m81_4/bb[6]_uq0 saout_m2_3v256x8m81_4/bb[7]_uq0
+ saout_m2_3v256x8m81_4/bb[5] saout_m2_3v256x8m81_4/bb[4]_uq0 saout_m2_3v256x8m81_4/bb[1]_uq0
+ saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_4/b[6] bb[10] ypass[2] WEN[1] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ b[12] men saout_m2_3v256x8m81_4/outbuf_oe_3v256x8m81_0/GWE b[10] ypass[0] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ b[9] bb[11] ypass[5] b[6] ypass[1] saout_m2_3v256x8m81_4/b[3] ypass[4] bb[8] saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ VDD_uq1 ypass[3] VSS ypass[7] ypass[6] VDD_uq0 VDD_uq4 VDD saout_m2_3v256x8m81
.ends

.subckt dcap_103_novia_3v256x8m81 w_n205_0# a_n30_42# a_n119_86#
X0 a_n119_86# a_n30_42# a_n119_86# w_n205_0# pfet_03v3 ad=0.4717p pd=3.01u as=0 ps=0 w=1.06u l=1.74u
.ends

.subckt lcol4_256_3v256x8m81 WL[20] WL[19] WL[18] WL[16] WL[14] WL[13] WL[12] WL[10]
+ WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[31] din[1] din[3] din[2]
+ q[1] q[2] q[3] pcb[2] pcb[3] pcb[0] pcb[1] WEN[3] WEN[2] WEN[1] WEN[0] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/outbuf_oe_3v256x8m81_0/GWE
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/q col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/q
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/GWEN col_256a_3v256x8m81_0/WL[6] col_256a_3v256x8m81_0/WL[8]
+ col_256a_3v256x8m81_0/WL[21] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/datain
+ WL[21] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/vdd_uq4 WL[22] WL[23] WL[24]
+ WL[25] WL[26] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/datain WL[27] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/datain
+ WL[28] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/q col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/q
+ col_256a_3v256x8m81_0/ypass[0] col_256a_3v256x8m81_0/ypass[1] col_256a_3v256x8m81_0/ypass[2]
+ col_256a_3v256x8m81_0/GWE col_256a_3v256x8m81_0/ypass[3] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/GWE
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/datain col_256a_3v256x8m81_0/ypass[4]
+ col_256a_3v256x8m81_0/men col_256a_3v256x8m81_0/WL[10] col_256a_3v256x8m81_0/ypass[5]
+ WL[11] col_256a_3v256x8m81_0/ypass[6] col_256a_3v256x8m81_0/ypass[7] col_256a_3v256x8m81_0/WL[12]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/GWE col_256a_3v256x8m81_0/VDD_uq5
+ WL[29] col_256a_3v256x8m81_0/WL[13] col_256a_3v256x8m81_0/VDD_uq3 col_256a_3v256x8m81_0/WL[14]
+ WL[30] col_256a_3v256x8m81_0/VDD_uq2 col_256a_3v256x8m81_0/WL[15] col_256a_3v256x8m81_0/VDD
+ WL[15] col_256a_3v256x8m81_0/VDD_uq1 col_256a_3v256x8m81_0/WL[17] col_256a_3v256x8m81_0/VDD_uq4
+ WL[17] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/GWE WL[0] VSUBS col_256a_3v256x8m81_0/WL[19]
+ col_256a_3v256x8m81_0/VDD_uq0 VDD
Xldummy_3v256x4_3v256x8m81_0 WL[5] VDD VSUBS col_256a_3v256x8m81_0/b[16] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ col_256a_3v256x8m81_0/b[16] VDD col_256a_3v256x8m81_0/bb[10] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ col_256a_3v256x8m81_0/WL[21] VDD WL[25] col_256a_3v256x8m81_0/b[10] col_256a_3v256x8m81_0/b[29]
+ VSUBS VSUBS col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[5] VDD col_256a_3v256x8m81_0/WL[6]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/b[3] VSUBS col_256a_3v256x8m81_0/bb[10]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/b[6] col_256a_3v256x8m81_0/b[10] WL[7]
+ WL[3] VDD VSUBS VSUBS col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ WL[23] VDD WL[22] VSUBS VSUBS col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[4] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/bb[2]
+ WL[4] VSUBS col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ col_256a_3v256x8m81_0/b[31] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ WL[9] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ VSUBS VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[1] col_256a_3v256x8m81_0/bb[24]
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[1] col_256a_3v256x8m81_0/bb[24] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ VDD col_256a_3v256x8m81_0/b[5] WL[21] WL[24] VSUBS VSUBS col_256a_3v256x8m81_0/bb[30]
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[6] WL[0] VSUBS VSUBS col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[7] col_256a_3v256x8m81_0/bb[6]
+ WL[11] VSUBS VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[2] col_256a_3v256x8m81_0/b[25]
+ VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[2] col_256a_3v256x8m81_0/b[25]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/bb[4] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ VDD VDD WL[19] WL[26] col_256a_3v256x8m81_0/b[31] VSUBS VSUBS col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/b[3] WL[2] VSUBS col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ col_256a_3v256x8m81_0/bb[11] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/b[6]
+ col_256a_3v256x8m81_0/WL[13] VSUBS VDD VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[3]
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[3] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ VDD VDD col_256a_3v256x8m81_0/bb[4] WL[17] VSUBS WL[28] VSUBS col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[7] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[4] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/bb[5]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ col_256a_3v256x8m81_0/WL[15] VSUBS VDD col_256a_3v256x8m81_0/b[29] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[5]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/b[3] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/b[6]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ VDD WL[15] VSUBS col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/b[12] VDD col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[5]
+ col_256a_3v256x8m81_0/WL[17] VSUBS VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[4] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[4]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/bb[2] VDD col_256a_3v256x8m81_0/WL[14]
+ VSUBS col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/b[6] VDD col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[5] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ VSUBS col_256a_3v256x8m81_0/WL[12] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ col_256a_3v256x8m81_0/bb[6] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ WL[30] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ VSUBS col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/b[3] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ WL[29] col_256a_3v256x8m81_0/bb[30] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/b[3]
+ VSUBS col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[6] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ col_256a_3v256x8m81_0/WL[10] VSUBS col_256a_3v256x8m81_0/bb[11] VDD col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/b[3] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ col_256a_3v256x8m81_0/b[5] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ VDD VDD col_256a_3v256x8m81_0/b[18] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ WL[27] col_256a_3v256x8m81_0/bb[8] VSUBS col_256a_3v256x8m81_0/b[18] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ col_256a_3v256x8m81_0/WL[8] VSUBS VDD col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/bb[4] col_256a_3v256x8m81_0/bb[8]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/bb[5] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ WL[1] col_256a_3v256x8m81_0/bb[17] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ col_256a_3v256x8m81_0/bb[17] VDD col_256a_3v256x8m81_0/b[9] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ VDD col_256a_3v256x8m81_0/WL[19] VSUBS col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[3]
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[3] VSUBS col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ col_256a_3v256x8m81_0/b[9] VDD col_256a_3v256x8m81_0/b[12] col_256a_3v256x8m81_0/bb[4]
+ ldummy_3v256x4_3v256x8m81
Xcol_256a_3v256x8m81_0 col_256a_3v256x8m81_0/ypass[0] col_256a_3v256x8m81_0/ypass[1]
+ col_256a_3v256x8m81_0/ypass[3] col_256a_3v256x8m81_0/ypass[4] col_256a_3v256x8m81_0/ypass[5]
+ col_256a_3v256x8m81_0/ypass[7] col_256a_3v256x8m81_0/VDD VSUBS WL[30] WL[29] WL[19]
+ WL[11] col_256a_3v256x8m81_0/WL[10] WL[7] WL[17] col_256a_3v256x8m81_0/WL[17] WL[15]
+ col_256a_3v256x8m81_0/WL[15] col_256a_3v256x8m81_0/WL[14] col_256a_3v256x8m81_0/WL[13]
+ WL[26] WL[25] col_256a_3v256x8m81_0/ypass[6] col_256a_3v256x8m81_0/ypass[2] col_256a_3v256x8m81_0/b[1]
+ col_256a_3v256x8m81_0/b[7] col_256a_3v256x8m81_0/b[10] col_256a_3v256x8m81_0/b[13]
+ col_256a_3v256x8m81_0/b[16] col_256a_3v256x8m81_0/b[22] col_256a_3v256x8m81_0/b[28]
+ col_256a_3v256x8m81_0/din[1] col_256a_3v256x8m81_0/din[3] col_256a_3v256x8m81_0/din[2]
+ col_256a_3v256x8m81_0/din[0] col_256a_3v256x8m81_0/q[0] col_256a_3v256x8m81_0/q[1]
+ col_256a_3v256x8m81_0/q[2] col_256a_3v256x8m81_0/q[3] col_256a_3v256x8m81_0/b[29]
+ col_256a_3v256x8m81_0/b[23] col_256a_3v256x8m81_0/b[20] col_256a_3v256x8m81_0/b[14]
+ col_256a_3v256x8m81_0/b[11] col_256a_3v256x8m81_0/b[8] col_256a_3v256x8m81_0/bb[0]
+ col_256a_3v256x8m81_0/bb[1] col_256a_3v256x8m81_0/bb[2] col_256a_3v256x8m81_0/bb[8]
+ col_256a_3v256x8m81_0/bb[9] col_256a_3v256x8m81_0/bb[11] col_256a_3v256x8m81_0/bb[12]
+ col_256a_3v256x8m81_0/bb[13] col_256a_3v256x8m81_0/bb[14] col_256a_3v256x8m81_0/bb[15]
+ col_256a_3v256x8m81_0/bb[19] col_256a_3v256x8m81_0/bb[21] col_256a_3v256x8m81_0/bb[22]
+ col_256a_3v256x8m81_0/bb[24] col_256a_3v256x8m81_0/bb[26] col_256a_3v256x8m81_0/bb[28]
+ col_256a_3v256x8m81_0/bb[29] col_256a_3v256x8m81_0/bb[30] col_256a_3v256x8m81_0/bb[31]
+ col_256a_3v256x8m81_0/b[30] col_256a_3v256x8m81_0/b[27] col_256a_3v256x8m81_0/b[0]
+ col_256a_3v256x8m81_0/b[3] col_256a_3v256x8m81_0/b[18] col_256a_3v256x8m81_0/pcb[0]
+ col_256a_3v256x8m81_0/pcb[1] col_256a_3v256x8m81_0/pcb[3] col_256a_3v256x8m81_0/pcb[2]
+ WEN[3] WEN[2] WEN[1] WEN[0] col_256a_3v256x8m81_0/VDD_uq5 col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/q
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/datain col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/GWEN
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/outbuf_oe_3v256x8m81_0/GWE WL[1] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/q WL[4] col_256a_3v256x8m81_0/men col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/vdd_uq4
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ col_256a_3v256x8m81_0/WL[21] VSUBS col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/datain
+ col_256a_3v256x8m81_0/b[9] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ WL[23] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/GWE col_256a_3v256x8m81_0/VDD_uq4
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[6] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ col_256a_3v256x8m81_0/b[25] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ WL[5] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ col_256a_3v256x8m81_0/VDD_uq1 col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/GWE col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ col_256a_3v256x8m81_0/WL[8] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[1] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[5]
+ WL[24] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/b[6] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[5]
+ WL[2] WL[27] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/b[3] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[3]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/q col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/q WL[21] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/b[3]
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/datain col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ col_256a_3v256x8m81_0/b[31] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/GWE col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ col_256a_3v256x8m81_0/VDD_uq3 col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/bb[2]
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/VDD_uq2 WL[9] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ col_256a_3v256x8m81_0/bb[4] col_256a_3v256x8m81_0/WL[12] col_256a_3v256x8m81_0/b[12]
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/bb[5] col_256a_3v256x8m81_0/GWE col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ WL[3] col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[4] WL[28] col_256a_3v256x8m81_0/b[5]
+ col_256a_3v256x8m81_0/WL[6] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/bb[4]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/datain col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/b[3]
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ col_256a_3v256x8m81_0/bb[17] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/b[6] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[4]
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_4/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/bb[2] col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_0/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ col_256a_3v256x8m81_0/saout_m2_3v256x8m81_3/b[3] col_256a_3v256x8m81_0/VDD_uq0 WL[22]
+ col_256a_3v256x8m81_0/saout_R_m2_3v256x8m81_1/bb[7] col_256a_3v256x8m81_0/bb[10]
+ VSUBS col_256a_3v256x8m81_0/WL[19] VDD WL[0] col_256a_3v256x8m81_0/bb[6] col_256a_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[0] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[1] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[2] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[3] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[4] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[5] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[6] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[7] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[8] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[9] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[10] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[11] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[12] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[13] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[14] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[15] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[16] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[17] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[18] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[19] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[20] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[21] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[22] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[23] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[24] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[25] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[26] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[27] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[28] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[29] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[30] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[31] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[32] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[33] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[34] VDD VSUBS VDD dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[35] VDD VSUBS VDD dcap_103_novia_3v256x8m81
.ends

.subckt rarray4_256_3v256x8m81 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8281#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13129#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_19189#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11203# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16765#
+ m3_n1397_8779# m3_n1397_13627# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n1397_3931#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1009#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# m3_n1397_19687# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n1397_18475#
+ m3_n1397_15553# m3_n1397_9991# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ m3_n1397_3433# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n1397_12415#
+ m3_n1397_2719# m3_n1397_14839# m3_n1397_17977# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_10705#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_247# m3_n1397_1507# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ m3_n1397_5143# m3_n1397_5857# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n1397_9493#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n1397_11917#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# m3_n1397_6355# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n1397_7567#
+ m3_n1397_7069# m3_n1397_16051# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
X018SRAM_cell1_2x_3v256x8m81_456 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_467 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_423 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_412 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_434 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_445 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_478 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_401 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_990 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_7 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_220 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_231 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_297 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_286 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_253 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_275 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_242 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_264 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_19 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_457 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_424 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_413 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_468 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_435 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_446 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_479 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_402 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_980 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_8 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_221 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_210 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_298 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_287 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_254 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_276 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_243 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_265 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_232 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1020 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_425 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_414 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_469 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_447 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_458 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_436 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_403 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_9 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_992 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_970 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_200 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_222 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_211 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1010 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_299 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_288 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_255 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_277 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_244 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_266 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_233 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_448 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_426 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_415 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_437 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_459 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_404 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_982 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_960 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_201 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_234 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_223 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1000 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_245 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1022 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_212 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_278 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_289 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_267 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_449 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_416 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_438 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_405 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_427 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_994 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_972 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1012 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_235 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_202 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_257 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_279 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_246 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_268 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_224 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_213 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_439 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_417 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_406 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_428 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_984 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_962 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1002 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_203 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_258 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_269 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_247 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_214 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_225 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_236 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_418 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_429 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_407 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_996 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_974 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_204 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_226 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1014 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_259 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_248 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_215 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_237 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_419 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_408 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_986 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_964 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_216 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_205 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_227 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_238 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1004 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_249 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_409 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_998 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_976 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_217 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_206 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_239 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_228 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1016 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_988 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_966 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1006 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_207 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_229 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_218 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_390 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_978 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1018 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_208 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_219 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_391 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_380 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_968 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_209 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1008 m3_n1397_18475# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_19189# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_18475#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_19189# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_392 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_370 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_381 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_371 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_393 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_360 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_382 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_190 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_394 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_350 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_372 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_361 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_383 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_191 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_180 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_395 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_351 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_362 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_340 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_384 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_373 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_192 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_181 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_170 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_330 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_341 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_396 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_352 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_374 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_363 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_385 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_193 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_182 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_160 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_171 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_512 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_397 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_353 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_320 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_375 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_386 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_364 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_342 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_331 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_194 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_183 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_161 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_172 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_150 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_354 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_310 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_343 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_321 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_332 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_398 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_376 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_387 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_365 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_184 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_195 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_162 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_173 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_140 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_151 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_333 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_300 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_399 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_344 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_311 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_377 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_388 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_366 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_322 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_355 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_196 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_185 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_163 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_174 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_130 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_141 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_152 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_90 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_334 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_301 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_345 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_389 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_378 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_367 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_323 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_312 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_356 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_120 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_197 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_186 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_164 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_175 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_131 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_142 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_153 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_91 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_80 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_335 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_302 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_379 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_346 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_368 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_324 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_313 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_357 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_198 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_187 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_165 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_176 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_132 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_143 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_121 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_110 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_154 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_92 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_70 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_81 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_303 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_347 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_336 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_369 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_325 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_314 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_358 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_188 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_199 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_166 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_177 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_144 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_111 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_100 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_133 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_122 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_155 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_93 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_60 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_82 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_71 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_304 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_348 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_326 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_337 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_315 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_359 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_167 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_189 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_178 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_112 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_134 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_123 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_156 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_145 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_101 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_50 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_94 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_61 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_72 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_83 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_305 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_994/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_327 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_349 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_338 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_316 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_168 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_179 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_124 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_135 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_157 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_113 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_146 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_102 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_40 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_51 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_95 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_62 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_73 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_84 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_328 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_306 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_339 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_317 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_114 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_103 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_125 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_169 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_158 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_136 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_147 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_41 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_52 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_30 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_96 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_63 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_74 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_85 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_329 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_307 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_318 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_115 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_137 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_159 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_148 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_104 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_126 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_42 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_53 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_20 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_31 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_64 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_75 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_86 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_97 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_319 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_308 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_457/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_116 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_138 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_127 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_149 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_82/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_105 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_43 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_10 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_54 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_21 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_32 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_65 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_87 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_98 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_76 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_309 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_139 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_106 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_128 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_117 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_470 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_44 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_11 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_55 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_22 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_33 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_99 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_88 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_98/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_66 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_77 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_118 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_96/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_129 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_107 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_471 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_460 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_290 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_45 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_12 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_34 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_23 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_56 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_67 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_78 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_89 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_108 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_119 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_99/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_472 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_461 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_998/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_450 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_280 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_291 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_46 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_46/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_13 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_35 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_24 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_57 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_68 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_79 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_81/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_109 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_65/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_451 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_440 m3_n1397_16051# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_16765# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_16051#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_16765# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_462 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_473 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_292 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_281 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_270 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_14 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_47 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_36 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_25 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_58 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_69 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_89/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_452 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_430 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_463 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_441 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_474 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_976/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_260 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_282 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_293 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_271 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_15 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_48 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_37 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_26 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_59 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_62/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_464 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_467/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_475 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_475/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_453 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_996/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_420 m3_n1397_17263# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_17977# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_17263#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_17977# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_431 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_442 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_4 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_261 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_283 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_250 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_294 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_272 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_49 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_38 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_27 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_16 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_476 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_454 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_421 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_465 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_410 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_443 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_432 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_5 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_9/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_262 m3_n1397_6355# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_7069# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_6355#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_7069# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_284 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_251 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_295 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_240 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_273 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_39 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_49/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_17 m3_n1397_1507# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_2221# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_1507#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_2221# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_28 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_477 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_477/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_455 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_422 m3_n1397_12415# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_13129# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_12415#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_13129# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_411 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_466 m3_n1397_9991# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_10705# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_9991#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_972/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_10705# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_433 m3_n1397_13627# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_14341# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_13627#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_14341# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_444 m3_n1397_14839# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_15553# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_14839#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_970/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_15553# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_400 m3_n1397_11203# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_11917# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_11203#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_11917# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_6 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_230 m3_n1397_8779# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_9493# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_8779#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_55/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_9493# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_296 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_992/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_263 m3_n1397_7567# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_8281# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_7567#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_966/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_8281# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_285 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_964/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_252 m3_n1397_2719# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_3433# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_2719#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_974/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_3433# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_241 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_968/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_274 m3_n1397_3931# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_4645# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_3931#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_978/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_4645# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_18 m3_n1397_247# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_1009# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_247#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_23/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_1009# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_29 m3_n1397_5143# VSUBS 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# VSUBS m3_n1397_5857# 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512#
+ 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n1397_5143#
+ 018SRAM_strap1_bndry_3v256x8m81_9/w_91_512# 018SRAM_cell1_2x_3v256x8m81_33/018SRAM_cell1_3v256x8m81_1/a_430_96#
+ m3_n1397_5857# VSUBS x018SRAM_cell1_2x_3v256x8m81
.ends

.subckt x018SRAM_cell1_dummy_R_3v256x8m81 m3_82_330# a_248_342# a_62_178# w_30_512#
+ a_430_96# a_110_96# a_192_298# VSUBS
X0 a_192_298# a_192_298# a_110_250# w_30_512# pfet_03v3 ad=0.1613p pd=1.39u as=0.1238p ps=1.44u w=0.28u l=0.28u
X1 a_248_342# a_192_298# a_110_250# VSUBS nfet_03v3 ad=0.171p pd=1.33u as=0.15665p ps=1.32u w=0.45u l=0.28u
X2 a_408_342# a_248_342# a_192_298# w_30_512# pfet_03v3 ad=0.1238p pd=1.44u as=0.1613p ps=1.39u w=0.28u l=0.28u
X3 a_408_342# a_248_342# a_248_342# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.171p ps=1.33u w=0.45u l=0.28u
X4 a_110_250# a_62_178# a_110_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
X5 a_408_342# a_62_178# a_430_96# VSUBS nfet_03v3 ad=0.15665p pd=1.32u as=0.1208p ps=1.42u w=0.28u l=0.36u
.ends

.subckt pmos_5p04310591302095_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.4251p pd=2.155u as=0.7194p ps=4.15u w=1.635u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.7194p pd=4.15u as=0.4251p ps=2.155u w=1.635u l=0.28u
.ends

.subckt nmos_5p04310591302098_3v256x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.1664p pd=1.16u as=0.2816p ps=2.16u w=0.64u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.2816p pd=2.16u as=0.1664p ps=1.16u w=0.64u l=0.28u
.ends

.subckt pmos_5p04310591302097_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=1.2909p pd=5.485u as=2.1846p ps=10.81u w=4.965u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=2.1846p pd=10.81u as=1.2909p ps=5.485u w=4.965u l=0.28u
.ends

.subckt ypass_gate_3v256x8m81_0 bb db ypass d pcb m3_0_2091# pmos_5p0431059130201_3v256x8m81_2/D
+ m3_0_2831# vss a_64_1295# m3_0_3056# pmos_5p0431059130201_3v256x8m81_0/D m3_0_3781#
+ m3_0_1632# m3_0_3536# b m3_0_3291# VSUBS m3_0_2331# vdd m3_0_2581# vdd_uq0
Xnmos_5p0431059130202_3v256x8m81_0 nmos_5p0431059130202_3v256x8m81_0/D a_64_1295#
+ a_64_1295# VSUBS VSUBS VSUBS nmos_5p0431059130202_3v256x8m81
Xpmos_5p0431059130201_3v256x8m81_0 pmos_5p0431059130201_3v256x8m81_0/D nmos_5p0431059130202_3v256x8m81_0/D
+ vdd_uq0 b pmos_5p0431059130201_3v256x8m81
Xpmos_5p0431059130201_3v256x8m81_1 b pcb vdd bb pmos_5p0431059130201_3v256x8m81
Xpmos_5p0431059130201_3v256x8m81_2 pmos_5p0431059130201_3v256x8m81_2/D nmos_5p0431059130202_3v256x8m81_0/D
+ vdd bb pmos_5p0431059130201_3v256x8m81
Xnmos_5p0431059130200_3v256x8m81_0 pmos_5p0431059130201_3v256x8m81_2/D a_64_1295#
+ bb VSUBS nmos_5p0431059130200_3v256x8m81
Xnmos_5p0431059130200_3v256x8m81_1 pmos_5p0431059130201_3v256x8m81_0/D a_64_1295#
+ b VSUBS nmos_5p0431059130200_3v256x8m81
X0 vdd pcb b vdd pfet_03v3 ad=0.94105p pd=4.37u as=0.51437p ps=2.24u w=1.595u l=0.28u
X1 bb pcb vdd vdd pfet_03v3 ad=0.51437p pd=2.24u as=1.13245p ps=4.61u w=1.595u l=0.28u
X2 nmos_5p0431059130202_3v256x8m81_0/D a_64_1295# vdd_uq0 vdd_uq0 pfet_03v3 ad=0.1946p pd=1.255u as=0.38225p ps=2.49u w=0.695u l=0.28u
X3 vdd_uq0 a_64_1295# nmos_5p0431059130202_3v256x8m81_0/D vdd_uq0 pfet_03v3 ad=0.50735p pd=2.85u as=0.1946p ps=1.255u w=0.695u l=0.28u
X4 b pcb vdd vdd pfet_03v3 ad=0.51437p pd=2.24u as=1.13245p ps=4.61u w=1.595u l=0.28u
X5 vdd pcb bb vdd pfet_03v3 ad=0.94105p pd=4.37u as=0.51437p ps=2.24u w=1.595u l=0.28u
.ends

.subckt nmos_5p04310591302096_3v256x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=1.0309p pd=4.485u as=1.7446p ps=8.81u w=3.965u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=1.7446p pd=8.81u as=1.0309p ps=4.485u w=3.965u l=0.28u
.ends

.subckt rdummy_3v256x4_3v256x8m81 018SRAM_cell1_dummy_3v256x8m81_62/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_23/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_33/w_30_512# ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_3v256x8m81_62/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_23/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ pmos_5p04310591302097_3v256x8m81_0/D m3_15667_n5798# 018SRAM_cell1_dummy_R_3v256x8m81_8/a_192_298#
+ 018SRAM_cell1_dummy_3v256x8m81_33/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_33/m2_134_89# 018SRAM_cell1_dummy_R_3v256x8m81_3/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_0/018SRAM_cell1_3v256x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_0/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_43/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_43/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_7/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_7/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89# 018SRAM_cell1_dummy_R_3v256x8m81_2/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/m3_82_330# w_15880_n13729#
+ 018SRAM_cell1_dummy_3v256x8m81_53/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_53/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_63/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_24/m2_346_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_0/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_63/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_24/m2_134_89# 018SRAM_cell1_dummy_R_3v256x8m81_10/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_10/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_6/a_192_298#
+ 018SRAM_cell1_dummy_3v256x8m81_34/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_34/m2_134_89# 018SRAM_cell1_dummy_R_3v256x8m81_40/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_0/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_0/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_44/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_44/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_30/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_8/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_30/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_8/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/w_30_512# 018SRAM_cell1_dummy_R_3v256x8m81_33/a_192_298#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89# m1_16100_n16182# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_54/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_54/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_40/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_40/a_248_342# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_dummy_3v256x8m81_64/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_25/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_64/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_25/m2_134_89# 018SRAM_cell1_dummy_R_3v256x8m81_11/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/w_30_512# 018SRAM_cell1_dummy_R_3v256x8m81_11/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_2/a_192_298# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_dummy_3v256x8m81_35/m2_346_89#
+ 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_35/m2_134_89#
+ ypass_gate_3v256x8m81_0_0/vss 018SRAM_cell1_dummy_R_3v256x8m81_38/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_45/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_45/m2_134_89# 018SRAM_cell1_dummy_R_3v256x8m81_9/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_9/a_248_342# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ ypass_gate_3v256x8m81_0_0/vdd 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_dummy_3v256x8m81_55/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_16/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_55/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_16/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/a_248_342# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_26/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_26/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_12/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v256x8m81_12/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_4/a_192_298#
+ 018SRAM_cell1_dummy_3v256x8m81_36/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_36/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_dummy_R_3v256x8m81_4/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_16/018SRAM_cell1_3v256x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_16/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_46/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_46/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/w_30_512# 018SRAM_cell1_dummy_R_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_17/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_56/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_56/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_17/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ m3_15667_n5552# 018SRAM_cell1_dummy_3v256x8m81_27/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v256x8m81_34/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_27/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/w_30_512# 018SRAM_cell1_dummy_R_3v256x8m81_13/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_13/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_7/a_192_298#
+ 018SRAM_cell1_dummy_3v256x8m81_37/m2_346_89# ypass_gate_3v256x8m81_0_0/vdd_uq0 018SRAM_cell1_dummy_3v256x8m81_37/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_16/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_16/018SRAM_cell1_3v256x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_65/a_192_298#
+ 018SRAM_cell1_dummy_3v256x8m81_47/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_47/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_33/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/w_30_512# ypass_gate_3v256x8m81_0_0/pmos_5p0431059130201_3v256x8m81_0/D
+ 018SRAM_cell1_dummy_R_3v256x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_33/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_57/m2_346_89#
+ m3_15667_n6510# 018SRAM_cell1_dummy_3v256x8m81_18/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89#
+ pmos_5p04310591302095_3v256x8m81_0/S 018SRAM_cell1_dummy_3v256x8m81_18/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_57/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_0/m3_82_330# 018SRAM_cell1_dummy_3v256x8m81_28/m2_346_89#
+ 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_39/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_28/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v256x8m81_14/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_14/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_5/a_192_298# 018SRAM_cell1_dummy_3v256x8m81_38/m2_346_89#
+ m3_15667_n6288# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_38/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_48/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_15/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_48/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_15/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_dummy_R_3v256x8m81_34/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_34/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_19/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_19/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_29/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_7/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_29/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_15/m3_82_330# m3_15698_n15942# 018SRAM_cell1_dummy_R_3v256x8m81_15/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_3/a_192_298# 018SRAM_cell1_dummy_3v256x8m81_39/m2_346_89#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_dummy_3v256x8m81_39/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_25/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_8/w_30_512# 018SRAM_cell1_dummy_R_3v256x8m81_25/a_248_342#
+ m3_15667_n7247# 018SRAM_cell1_dummy_R_3v256x8m81_40/a_192_298# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_dummy_3v256x8m81_49/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_15/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_49/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_15/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_2/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_35/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_2/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_35/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_38/a_192_298# 018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_59/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_dummy_3v256x8m81_59/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v256x8m81_16/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_2/018SRAM_cell1_3v256x8m81_0/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_16/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_2/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_65/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_26/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_65/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_26/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_34/a_192_298#
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_3/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_3/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_14/018SRAM_cell1_3v256x8m81_0/m3_82_330# 018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ m3_15645_n13711# 018SRAM_cell1_dummy_R_3v256x8m81_39/a_192_298# 018SRAM_cell1_2x_3v256x8m81_14/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_20/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_20/m2_134_89# 018SRAM_cell1_dummy_R_3v256x8m81_17/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_2/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_17/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_2/018SRAM_cell1_3v256x8m81_1/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_30/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_30/m2_134_89# 018SRAM_cell1_dummy_R_3v256x8m81_27/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_65/w_30_512# 018SRAM_cell1_dummy_R_3v256x8m81_27/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_40/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_40/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_4/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ 018SRAM_cell1_dummy_R_3v256x8m81_4/a_248_342# 018SRAM_cell1_2x_3v256x8m81_14/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_14/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_3v256x8m81_50/m2_346_89# 018SRAM_cell1_dummy_R_3v256x8m81_5/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_50/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_3v256x8m81_21/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_60/m2_346_89#
+ 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_6/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_60/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_21/m2_134_89#
+ 018SRAM_cell1_dummy_R_3v256x8m81_18/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_18/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_dummy_R_3v256x8m81_0/a_192_298#
+ 018SRAM_cell1_dummy_3v256x8m81_31/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_1/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ m3_15667_n6043# 018SRAM_cell1_dummy_3v256x8m81_31/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_1/018SRAM_cell1_3v256x8m81_0/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_28/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_28/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_dummy_3v256x8m81_41/m2_346_89#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_0/m3_82_330# 018SRAM_cell1_dummy_3v256x8m81_41/m2_134_89#
+ m2_16574_19394# 018SRAM_cell1_dummy_R_3v256x8m81_38/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_5/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_5/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_38/a_248_342# 018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_51/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_51/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_61/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_22/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_22/m2_134_89# 018SRAM_cell1_dummy_3v256x8m81_61/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/m3_82_330# a_n547_178#
+ 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_1/a_192_298#
+ 018SRAM_cell1_dummy_3v256x8m81_32/m2_346_89# 018SRAM_cell1_2x_3v256x8m81_1/018SRAM_cell1_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_dummy_3v256x8m81_32/m2_134_89# 018SRAM_cell1_2x_3v256x8m81_1/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_29/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_29/a_248_342#
+ m3_15667_n7002# pmos_5p04310591302097_3v256x8m81_0/S 018SRAM_cell1_dummy_3v256x8m81_42/m2_346_89#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# 018SRAM_cell1_dummy_3v256x8m81_42/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_dummy_R_3v256x8m81_39/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_6/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_dummy_R_3v256x8m81_39/a_248_342# 018SRAM_cell1_dummy_R_3v256x8m81_6/a_248_342#
+ m2_16574_21# 018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_52/m2_346_89#
+ m3_n631_83# 018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89# 018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89#
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/a_248_592# ypass_gate_3v256x8m81_0_0/pcb
+ 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/w_30_512# VSUBS 018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89#
+ 018SRAM_cell1_dummy_3v256x8m81_52/m2_134_89# m3_15667_n6752#
X018SRAM_cell1_2x_3v256x8m81_7 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n631_83# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n631_83# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_5 018SRAM_cell1_dummy_R_3v256x8m81_5/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_5/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_5/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_5/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_19 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n631_83# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n631_83# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_54 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_54/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_54/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_43 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_43/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_43/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_32 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_32/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_32/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_21 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_21/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_21/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_10 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_10/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_10/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_25 018SRAM_cell1_dummy_R_3v256x8m81_25/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_25/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_33/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_33/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_14 018SRAM_cell1_dummy_R_3v256x8m81_14/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_14/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_2/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_2/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_6 018SRAM_cell1_dummy_R_3v256x8m81_6/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_6/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_6/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_6/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_8 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n631_83# 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n631_83# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_55 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_55/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_55/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_44 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_44/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_44/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_33 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_33/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_33/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_22 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_22/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_22/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_11 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_11/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_11/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_26 018SRAM_cell1_dummy_R_3v256x8m81_26/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_26/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_65/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_65/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_15 018SRAM_cell1_dummy_R_3v256x8m81_15/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_15/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_4/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_4/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_7 018SRAM_cell1_dummy_R_3v256x8m81_7/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_7/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_7/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_7/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
Xpmos_5p04310591302095_3v256x8m81_0 pmos_5p04310591302095_3v256x8m81_0/D ypass_gate_3v256x8m81_0_0/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_0_0/pmos_5p0431059130201_3v256x8m81_0/D pmos_5p04310591302095_3v256x8m81_0/S
+ pmos_5p04310591302095_3v256x8m81_0/S pmos_5p04310591302095_3v256x8m81_0/S pmos_5p04310591302095_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_56 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_56/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_56/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_45 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_45/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_45/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_34 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_34/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_34/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_23 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_23/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_23/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_12 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_12/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_12/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_27 018SRAM_cell1_dummy_R_3v256x8m81_27/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_27/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_38/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_38/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_38 018SRAM_cell1_dummy_R_3v256x8m81_38/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_38/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_38/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_38/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_16 018SRAM_cell1_dummy_R_3v256x8m81_16/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_16/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_7/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_7/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_8 018SRAM_cell1_dummy_R_3v256x8m81_8/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_8/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_8/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_8/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_57 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_57/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_57/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_46 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_46/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_46/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_35 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_35/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_35/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_24 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_24/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_24/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_13 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_13/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_13/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_28 018SRAM_cell1_dummy_R_3v256x8m81_28/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_28/a_248_342# m2_16574_19394# 018SRAM_cell1_dummy_R_3v256x8m81_40/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_40/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_39 018SRAM_cell1_dummy_R_3v256x8m81_39/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_39/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_39/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_39/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_17 018SRAM_cell1_dummy_R_3v256x8m81_17/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_17/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_5/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_5/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_9 018SRAM_cell1_dummy_R_3v256x8m81_9/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_9/a_248_342# m2_16574_21# 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_47 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_47/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_47/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_36 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_36/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_36/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_25 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_25/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_25/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_14 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_14/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_14/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_29 018SRAM_cell1_dummy_R_3v256x8m81_29/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_29/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_34/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_34/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_18 018SRAM_cell1_dummy_R_3v256x8m81_18/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_18/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_3/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_3/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_59 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_59/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_59/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_48 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_48/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_48/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_37 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_37/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_37/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_26 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_26/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_26/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_15 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_15/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_15/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_19 a_n547_178# VSUBS m2_16574_21# 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_49 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_49/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_49/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_38 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_38/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_38/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_27 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_27/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_27/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_16 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_16/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_16/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_39 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_39/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_39/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_28 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_28/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_28/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_17 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_17/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_17/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
Xnmos_5p04310591302098_3v256x8m81_0 pmos_5p04310591302095_3v256x8m81_0/D ypass_gate_3v256x8m81_0_0/pmos_5p0431059130201_3v256x8m81_0/D
+ ypass_gate_3v256x8m81_0_0/pmos_5p0431059130201_3v256x8m81_0/D VSUBS VSUBS VSUBS
+ nmos_5p04310591302098_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_29 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_29/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_29/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_18 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_18/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_18/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_19 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_19/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_19/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_0 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_0/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_0/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_3v256x8m81_0 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ a_n547_178# 018SRAM_cell1_3v256x8m81_0/w_30_512# 018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# VSUBS x018SRAM_cell1_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_1 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_1/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_1/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
Xpmos_5p04310591302097_3v256x8m81_0 pmos_5p04310591302097_3v256x8m81_0/D pmos_5p04310591302095_3v256x8m81_0/D
+ pmos_5p04310591302095_3v256x8m81_0/D w_15880_n13729# pmos_5p04310591302097_3v256x8m81_0/S
+ pmos_5p04310591302097_3v256x8m81_0/S pmos_5p04310591302097_3v256x8m81
X018SRAM_cell1_3v256x8m81_1 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ m3_n631_83# 018SRAM_cell1_3v256x8m81_1/w_30_512# 018SRAM_cell1_3v256x8m81_1/a_430_96#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# VSUBS x018SRAM_cell1_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_2 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_2/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_2/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_3 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_3/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_3/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
Xypass_gate_3v256x8m81_0_0 ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/db
+ ypass_gate_3v256x8m81_0_0/ypass ypass_gate_3v256x8m81_0_0/d ypass_gate_3v256x8m81_0_0/pcb
+ m3_15667_n7247# ypass_gate_3v256x8m81_0_0/bb m3_15667_n6510# ypass_gate_3v256x8m81_0_0/vss
+ ypass_gate_3v256x8m81_0_0/vdd_uq0 m3_15667_n6288# ypass_gate_3v256x8m81_0_0/pmos_5p0431059130201_3v256x8m81_0/D
+ m3_15667_n5552# ypass_gate_3v256x8m81_0_0/vdd_uq0 m3_15667_n5798# ypass_gate_3v256x8m81_0_0/b
+ m3_15667_n6043# VSUBS m3_15667_n7002# ypass_gate_3v256x8m81_0_0/vdd m3_15667_n6752#
+ ypass_gate_3v256x8m81_0_0/vdd_uq0 ypass_gate_3v256x8m81_0
X018SRAM_cell1_dummy_3v256x8m81_4 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_4/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_4/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_5 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_5/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_5/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_6 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_6/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_6/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_7 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_7/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_7/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_8 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_8/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_8/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_9 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_9/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_9/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_31 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n631_83# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n631_83# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_0 018SRAM_cell1_2x_3v256x8m81_0/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_0/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_0/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_0/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n631_83# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n631_83# VSUBS x018SRAM_cell1_2x_3v256x8m81
Xnmos_5p04310591302096_3v256x8m81_0 pmos_5p04310591302097_3v256x8m81_0/D pmos_5p04310591302095_3v256x8m81_0/D
+ pmos_5p04310591302095_3v256x8m81_0/D VSUBS VSUBS VSUBS nmos_5p04310591302096_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_40 018SRAM_cell1_dummy_R_3v256x8m81_40/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_40/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_40/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_40/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_1 018SRAM_cell1_2x_3v256x8m81_1/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_1/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_1/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_1/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n631_83# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n631_83# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_52 m2_16574_19394# VSUBS m2_16574_19394# 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_30 018SRAM_cell1_dummy_R_3v256x8m81_30/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_30/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_39/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_39/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_2 018SRAM_cell1_2x_3v256x8m81_2/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_2/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_2/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_2/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n631_83# 018SRAM_cell1_2x_3v256x8m81_7/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n631_83# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_0 018SRAM_cell1_dummy_R_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_0/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_0/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_0/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_60 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_60/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_60/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_14 018SRAM_cell1_2x_3v256x8m81_14/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_14/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_14/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_14/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n631_83# 018SRAM_cell1_2x_3v256x8m81_31/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n631_83# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_3 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_3/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n631_83# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n631_83# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_1 018SRAM_cell1_dummy_R_3v256x8m81_1/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_1/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_1/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_1/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_15 018SRAM_cell1_2x_3v256x8m81_15/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_15/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_15/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_15/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n631_83# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n631_83# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_61 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_61/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_61/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_50 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_50/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_50/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_65 018SRAM_cell1_dummy_R_3v256x8m81_65/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_65/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_65/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_65/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_10 018SRAM_cell1_dummy_R_3v256x8m81_10/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_10/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_0/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_0/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_4 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n631_83# 018SRAM_cell1_2x_3v256x8m81_4/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n631_83# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_2 018SRAM_cell1_dummy_R_3v256x8m81_2/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_2/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_2/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_2/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_62 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_62/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_62/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_51 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_51/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_51/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_40 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_40/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_40/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_16 018SRAM_cell1_2x_3v256x8m81_16/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_16/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_16/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_16/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n631_83# 018SRAM_cell1_2x_3v256x8m81_19/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n631_83# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_33 018SRAM_cell1_dummy_R_3v256x8m81_33/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_33/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_33/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_33/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_11 018SRAM_cell1_dummy_R_3v256x8m81_11/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_11/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_1/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_1/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_5 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n631_83# 018SRAM_cell1_2x_3v256x8m81_5/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n631_83# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_3 018SRAM_cell1_dummy_R_3v256x8m81_3/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_3/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_3/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_3/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_17 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n631_83# 018SRAM_cell1_2x_3v256x8m81_17/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n631_83# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_63 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_63/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_63/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_52 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_52/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_52/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_41 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_41/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_41/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_30 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_30/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_30/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_34 018SRAM_cell1_dummy_R_3v256x8m81_34/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_34/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_34/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_34/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_12 018SRAM_cell1_dummy_R_3v256x8m81_12/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_12/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_8/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_8/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_4 018SRAM_cell1_dummy_R_3v256x8m81_4/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_4/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_4/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_4/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_6 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/a_248_592# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_2x_3v256x8m81_6/018SRAM_cell1_3v256x8m81_1/a_248_592#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n631_83# 018SRAM_cell1_2x_3v256x8m81_8/018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n631_83# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_64 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_64/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_64/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_53 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_53/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_53/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_42 m2_16574_19394# VSUBS 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/w_30_512# m2_16574_19394# 018SRAM_cell1_dummy_3v256x8m81_42/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_42/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_2x_3v256x8m81_18 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/m3_82_330#
+ 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/a_248_342# 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/a_248_592# 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_1/a_248_342#
+ 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_1/m3_82_330# 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_110_96# m3_n631_83# 018SRAM_cell1_2x_3v256x8m81_18/018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_1/a_430_96# m3_n631_83# VSUBS x018SRAM_cell1_2x_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_31 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_31/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_31/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_3v256x8m81_20 a_n547_178# VSUBS 018SRAM_cell1_3v256x8m81_0/w_30_512#
+ 018SRAM_cell1_3v256x8m81_0/w_30_512# a_n547_178# 018SRAM_cell1_dummy_3v256x8m81_20/m2_346_89#
+ 018SRAM_cell1_dummy_3v256x8m81_20/m2_134_89# VSUBS x018SRAM_cell1_dummy_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_35 018SRAM_cell1_dummy_R_3v256x8m81_35/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_35/a_248_342# m2_16574_19394# 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_3v256x8m81_1/w_30_512#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
X018SRAM_cell1_dummy_R_3v256x8m81_13 018SRAM_cell1_dummy_R_3v256x8m81_13/m3_82_330#
+ 018SRAM_cell1_dummy_R_3v256x8m81_13/a_248_342# m2_16574_21# 018SRAM_cell1_dummy_R_3v256x8m81_6/w_30_512#
+ ypass_gate_3v256x8m81_0_0/bb ypass_gate_3v256x8m81_0_0/b 018SRAM_cell1_dummy_R_3v256x8m81_6/a_192_298#
+ VSUBS x018SRAM_cell1_dummy_R_3v256x8m81
.ends

.subckt rcol4_256_3v256x8m81 WL[29] WL[20] WL[27] WL[30] WL[18] WL[15] WL[31] WL[14]
+ WL[16] WL[26] WL[19] WL[28] WL[12] WL[8] WL[5] WL[10] WL[13] WL[6] tblhl GWE WL[11]
+ din[7] q[5] q[6] q[7] din[5] din[6] q[4] pcb[6] pcb[7] pcb[4] WEN[4] WEN[7] pcb[5]
+ WEN[5] WEN[6] rarray4_256_3v256x8m81_0/m3_n1397_10705# rdummy_3v256x4_3v256x8m81_0/ypass_gate_3v256x8m81_0_0/pcb
+ rarray4_256_3v256x8m81_0/m3_n1397_8779# rarray4_256_3v256x8m81_0/m3_n1397_8281#
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass saout_m2_3v256x8m81_2/datain
+ saout_m2_3v256x8m81_3/din_3v256x8m81_0/men saout_R_m2_3v256x8m81_1/datain saout_m2_3v256x8m81_2/q
+ rarray4_256_3v256x8m81_0/m3_n1397_13129# saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ rarray4_256_3v256x8m81_0/m3_n1397_11917# rarray4_256_3v256x8m81_0/m3_n1397_9493#
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass saout_R_m2_3v256x8m81_1/sa_3v256x8m81_0/pcb
+ rdummy_3v256x4_3v256x8m81_0/m2_16574_21# saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass
+ rarray4_256_3v256x8m81_0/m3_n1397_5143# WL[21] WL[7] rarray4_256_3v256x8m81_0/m3_n1397_3931#
+ WL[1] WL[0] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass
+ rarray4_256_3v256x8m81_0/m3_n1397_19687# saout_m2_3v256x8m81_3/VDD_uq0 rarray4_256_3v256x8m81_0/m3_n1397_6355#
+ saout_m2_3v256x8m81_3/vdd_uq0 WL[9] WL[23] WL[22] saout_m2_3v256x8m81_3/ypass[7]
+ saout_R_m2_3v256x8m81_1/q saout_m2_3v256x8m81_3/q WL[2] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass
+ saout_m2_3v256x8m81_3/vdd saout_m2_3v256x8m81_3/vdd_uq3 saout_R_m2_3v256x8m81_3/q
+ saout_R_m2_3v256x8m81_3/datain rarray4_256_3v256x8m81_0/m3_n1397_7567# WL[25] saout_R_m2_3v256x8m81_3/vdd
+ saout_m2_3v256x8m81_3/GWEN saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass
+ WL[24] saout_m2_3v256x8m81_3/vdd_uq2 saout_m2_3v256x8m81_3/datain WL[4] WL[3] WL[17]
+ saout_m2_3v256x8m81_3/VDD VSS saout_R_m2_3v256x8m81_3/b[7]
Xrarray4_256_3v256x8m81_0 saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b rarray4_256_3v256x8m81_0/m3_n1397_8281#
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_3/bb[3] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ rarray4_256_3v256x8m81_0/m3_n1397_13129# saout_R_m2_3v256x8m81_3/b[6] saout_m2_3v256x8m81_2/bb[5]
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b WL[30] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_m2_3v256x8m81_2/b[4] saout_R_m2_3v256x8m81_3/bb[2] saout_m2_3v256x8m81_3/b[4]
+ saout_m2_3v256x8m81_2/bb[3] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ WL[17] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb saout_R_m2_3v256x8m81_1/b[3]
+ saout_R_m2_3v256x8m81_3/bb[5] saout_m2_3v256x8m81_3/b[3] WL[26] rarray4_256_3v256x8m81_0/m3_n1397_8779#
+ WL[21] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ rarray4_256_3v256x8m81_0/m3_n1397_3931# saout_R_m2_3v256x8m81_1/b[6] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b WL[1] saout_R_m2_3v256x8m81_1/bb[7]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ WL[3] rarray4_256_3v256x8m81_0/m3_n1397_19687# saout_m2_3v256x8m81_3/bb[5] saout_R_m2_3v256x8m81_3/b[3]
+ WL[29] WL[24] WL[15] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ WL[5] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ saout_m2_3v256x8m81_2/b[3] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_m2_3v256x8m81_3/bb[2]
+ saout_R_m2_3v256x8m81_3/bb[4] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ WL[19] WL[4] WL[23] WL[28] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb rarray4_256_3v256x8m81_0/m3_n1397_10705#
+ saout_m2_3v256x8m81_3/b[1] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_R_m2_3v256x8m81_3/bb[7] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ WL[0] WL[2] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_R_m2_3v256x8m81_1/bb[5] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ WL[22] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b rarray4_256_3v256x8m81_0/m3_n1397_5143#
+ WL[9] saout_m2_3v256x8m81_2/b[1] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ rarray4_256_3v256x8m81_0/m3_n1397_9493# saout_R_m2_3v256x8m81_1/bb[2] rarray4_256_3v256x8m81_0/m3_n1397_11917#
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb WL[27] saout_m2_3v256x8m81_3/b[6]
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb WL[7] rarray4_256_3v256x8m81_0/m3_n1397_6355#
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_2/b[6] saout_R_m2_3v256x8m81_1/bb[4] rarray4_256_3v256x8m81_0/m3_n1397_7567#
+ WL[11] WL[25] saout_m2_3v256x8m81_2/bb[2] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ VSS saout_R_m2_3v256x8m81_3/b[7] rarray4_256_3v256x8m81
Xrdummy_3v256x4_3v256x8m81_0 saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb saout_R_m2_3v256x8m81_3/b[7]
+ rdummy_3v256x4_3v256x8m81_0/ypass_gate_3v256x8m81_0_0/b saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_3/b[7] WL[30] VSS tblhl saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/bb[5] saout_R_m2_3v256x8m81_3/b[7]
+ rarray4_256_3v256x8m81_0/m3_n1397_7567# VSS saout_R_m2_3v256x8m81_3/bb[4] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ rarray4_256_3v256x8m81_0/m3_n1397_8779# VSS saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_3/b[7] rarray4_256_3v256x8m81_0/m3_n1397_8779# saout_m2_3v256x8m81_3/vdd
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb saout_R_m2_3v256x8m81_1/bb[7]
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b VSS saout_m2_3v256x8m81_2/b[4]
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_3/b[1] saout_R_m2_3v256x8m81_3/b[7] saout_R_m2_3v256x8m81_1/bb[7]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb WL[5] VSS saout_R_m2_3v256x8m81_3/b[7]
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb WL[25] VSS
+ saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/b[4] saout_R_m2_3v256x8m81_3/b[7]
+ rarray4_256_3v256x8m81_0/m3_n1397_8281# VSS saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ saout_R_m2_3v256x8m81_3/bb[5] WL[25] rarray4_256_3v256x8m81_0/m3_n1397_7567# VSS
+ VSS saout_R_m2_3v256x8m81_3/b[7] saout_R_m2_3v256x8m81_3/b[7] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ tblhl rarray4_256_3v256x8m81_0/m3_n1397_9493# saout_m2_3v256x8m81_2/b[3] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ saout_R_m2_3v256x8m81_1/b[6] VSS saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_m2_3v256x8m81_2/bb[3] WL[28] WL[17] VSS VSS saout_R_m2_3v256x8m81_3/b[7] saout_R_m2_3v256x8m81_1/bb[2]
+ saout_m2_3v256x8m81_3/bb[2] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b WL[7] saout_R_m2_3v256x8m81_3/b[7]
+ VSS saout_R_m2_3v256x8m81_3/b[7] saout_R_m2_3v256x8m81_3/b[7] WL[26] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ VSS saout_m2_3v256x8m81_3/b[6] VSS saout_R_m2_3v256x8m81_3/b[7] saout_R_m2_3v256x8m81_3/b[3]
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb WL[0] VSS
+ saout_R_m2_3v256x8m81_3/b[7] saout_R_m2_3v256x8m81_3/b[7] saout_R_m2_3v256x8m81_3/b[7]
+ saout_m2_3v256x8m81_2/bb[2] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_R_m2_3v256x8m81_3/b[6]
+ rarray4_256_3v256x8m81_0/m3_n1397_6355# rarray4_256_3v256x8m81_0/m3_n1397_11917#
+ VSS VSS saout_m2_3v256x8m81_3/b[3] saout_m2_3v256x8m81_3/bb[3] WL[11] saout_R_m2_3v256x8m81_3/b[7]
+ VSS saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb saout_R_m2_3v256x8m81_3/b[7]
+ saout_R_m2_3v256x8m81_3/b[7] WL[23] VSS saout_R_m2_3v256x8m81_3/bb[2] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_R_m2_3v256x8m81_3/b[7] saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_3/bb[4] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ saout_R_m2_3v256x8m81_1/bb[5] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ WL[11] VSS saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b saout_R_m2_3v256x8m81_3/b[7]
+ saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/bb[5] saout_R_m2_3v256x8m81_3/b[7]
+ rarray4_256_3v256x8m81_0/m3_n1397_9493# VSS saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/b[1]
+ saout_m2_3v256x8m81_3/vdd_uq0 saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_R_m2_3v256x8m81_3/b[7] WL[24] VSS saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ rarray4_256_3v256x8m81_0/m3_n1397_3931# WL[22] saout_R_m2_3v256x8m81_3/b[7] rdummy_3v256x4_3v256x8m81_0/ypass_gate_3v256x8m81_0_0/b
+ VSS VSS saout_m2_3v256x8m81_2/b[1] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb saout_m2_3v256x8m81_3/vdd_uq3
+ saout_R_m2_3v256x8m81_3/bb[5] saout_R_m2_3v256x8m81_1/b[6] saout_R_m2_3v256x8m81_3/b[7]
+ WL[15] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb VSS
+ saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/b[4] saout_R_m2_3v256x8m81_3/b[7]
+ WL[3] VSS saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/bb[2] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass
+ WL[0] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b VSS saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ WL[27] saout_m2_3v256x8m81_2/bb[5] VSS rarray4_256_3v256x8m81_0/m3_n1397_5143# saout_R_m2_3v256x8m81_3/b[7]
+ WL[26] VSS VSS saout_m2_3v256x8m81_2/bb[2] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ saout_R_m2_3v256x8m81_3/b[3] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ rarray4_256_3v256x8m81_0/m3_n1397_10705# saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ VSS saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/b[6] WL[9] VSS VSS saout_R_m2_3v256x8m81_3/b[7]
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b WL[1] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ VSS WL[23] saout_R_m2_3v256x8m81_3/b[7] VSS saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass
+ saout_R_m2_3v256x8m81_3/b[7] saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_2/b[1]
+ WL[28] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb VSS
+ WL[4] WL[30] VSS VSS saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_2/b[3] saout_R_m2_3v256x8m81_1/b[3]
+ saout_m2_3v256x8m81_2/bb[3] saout_R_m2_3v256x8m81_3/b[7] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ saout_R_m2_3v256x8m81_3/b[7] rarray4_256_3v256x8m81_0/m3_n1397_8281# rarray4_256_3v256x8m81_0/m3_n1397_5143#
+ VSS VSS rarray4_256_3v256x8m81_0/m3_n1397_11917# WL[19] VSS VSS saout_R_m2_3v256x8m81_3/b[7]
+ rarray4_256_3v256x8m81_0/m3_n1397_3931# VSS WL[2] VSS WL[19] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_m2_3v256x8m81_3/vdd saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_1/bb[4]
+ saout_m2_3v256x8m81_2/bb[5] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b
+ WL[21] saout_R_m2_3v256x8m81_3/bb[2] VSS saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ rarray4_256_3v256x8m81_0/m3_n1397_10705# WL[9] VSS VSS saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb WL[21] saout_R_m2_3v256x8m81_3/b[7]
+ VSS WL[7] VSS saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_3/bb[7] rarray4_256_3v256x8m81_0/m3_n1397_6355# saout_R_m2_3v256x8m81_3/b[7]
+ VSS rarray4_256_3v256x8m81_0/m3_n1397_13129# saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb
+ VSS saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b saout_R_m2_3v256x8m81_3/b[7]
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_m2_3v256x8m81_2/b[4]
+ saout_R_m2_3v256x8m81_1/bb[5] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ saout_R_m2_3v256x8m81_3/b[7] WL[22] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b VSS saout_R_m2_3v256x8m81_3/b[7]
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ WL[1] VSS saout_R_m2_3v256x8m81_3/b[7] saout_R_m2_3v256x8m81_3/b[7] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ WL[4] saout_m2_3v256x8m81_3/ypass[7] saout_R_m2_3v256x8m81_3/bb[7] VSS WL[29] VSS
+ saout_R_m2_3v256x8m81_3/b[7] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ WL[2] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b rarray4_256_3v256x8m81_0/m3_n1397_19687#
+ rarray4_256_3v256x8m81_0/m3_n1397_13129# WL[17] VSS VSS VSS saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_R_m2_3v256x8m81_1/b[3] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_m2_3v256x8m81_2/b[6] saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_2/b[6]
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb saout_R_m2_3v256x8m81_1/bb[4]
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b WL[29] VSS
+ VSS saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/b[3] WL[5] saout_R_m2_3v256x8m81_3/b[7]
+ saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/bb[3] VSS WL[27] VSS saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass
+ saout_m2_3v256x8m81_3/vdd saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_R_m2_3v256x8m81_3/b[7] saout_R_m2_3v256x8m81_3/b[6] WL[3] WL[24] WL[15] VSS
+ VSS VSS rdummy_3v256x4_3v256x8m81_0/m2_16574_21# saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb VSS saout_R_m2_3v256x8m81_1/bb[2]
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb saout_R_m2_3v256x8m81_3/b[7]
+ rdummy_3v256x4_3v256x8m81_0/ypass_gate_3v256x8m81_0_0/pcb saout_R_m2_3v256x8m81_3/b[7]
+ VSS saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass rdummy_3v256x4_3v256x8m81
Xsaout_R_m2_3v256x8m81_1 saout_R_m2_3v256x8m81_1/ypass[2] saout_R_m2_3v256x8m81_1/ypass[3]
+ saout_R_m2_3v256x8m81_1/ypass[4] saout_R_m2_3v256x8m81_1/ypass[5] saout_R_m2_3v256x8m81_1/ypass[6]
+ saout_m2_3v256x8m81_3/GWEN saout_R_m2_3v256x8m81_1/datain saout_R_m2_3v256x8m81_1/b[5]
+ saout_R_m2_3v256x8m81_1/b[4] saout_R_m2_3v256x8m81_1/b[2] saout_R_m2_3v256x8m81_1/b[1]
+ saout_R_m2_3v256x8m81_1/b[0] saout_R_m2_3v256x8m81_1/bb[6] saout_R_m2_3v256x8m81_1/q
+ saout_R_m2_3v256x8m81_1/bb[3] saout_R_m2_3v256x8m81_1/bb[0] saout_R_m2_3v256x8m81_1/bb[1]
+ saout_R_m2_3v256x8m81_1/pcb saout_R_m2_3v256x8m81_1/vss_uq6 saout_m2_3v256x8m81_3/vdd_uq2
+ saout_R_m2_3v256x8m81_1/vdd_uq2 saout_R_m2_3v256x8m81_1/vdd_uq4 saout_R_m2_3v256x8m81_1/vdd_uq6
+ saout_R_m2_3v256x8m81_1/pcb_uq0 saout_R_m2_3v256x8m81_1/datain_uq0 saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_1/bb[5] saout_R_m2_3v256x8m81_1/sa_3v256x8m81_0/pcb saout_R_m2_3v256x8m81_1/sa_3v256x8m81_0/d
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b GWE saout_R_m2_3v256x8m81_1/bb[2]
+ WEN[4] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb saout_R_m2_3v256x8m81_1/b[3]
+ saout_m2_3v256x8m81_3/ypass[7] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass saout_R_m2_3v256x8m81_1/b[6]
+ saout_R_m2_3v256x8m81_1/bb[4] saout_R_m2_3v256x8m81_3/vdd saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass
+ saout_m2_3v256x8m81_3/din_3v256x8m81_0/men saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass
+ saout_R_m2_3v256x8m81_1/bb[7] saout_R_m2_3v256x8m81_1/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ saout_m2_3v256x8m81_3/vdd saout_m2_3v256x8m81_3/vdd_uq0 saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass
+ VSS saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass saout_m2_3v256x8m81_3/VDD
+ saout_m2_3v256x8m81_3/vdd_uq3 saout_m2_3v256x8m81_3/VDD_uq0 saout_R_m2_3v256x8m81
Xsaout_R_m2_3v256x8m81_3 saout_R_m2_3v256x8m81_3/ypass[2] saout_R_m2_3v256x8m81_3/ypass[3]
+ saout_R_m2_3v256x8m81_3/ypass[4] saout_R_m2_3v256x8m81_3/ypass[5] saout_R_m2_3v256x8m81_3/ypass[6]
+ saout_m2_3v256x8m81_3/GWEN saout_R_m2_3v256x8m81_3/datain saout_R_m2_3v256x8m81_3/b[5]
+ saout_R_m2_3v256x8m81_3/b[4] saout_R_m2_3v256x8m81_3/b[2] saout_R_m2_3v256x8m81_3/b[1]
+ saout_R_m2_3v256x8m81_3/b[0] saout_R_m2_3v256x8m81_3/bb[6] saout_R_m2_3v256x8m81_3/q
+ saout_R_m2_3v256x8m81_3/bb[3] saout_R_m2_3v256x8m81_3/bb[0] saout_R_m2_3v256x8m81_3/bb[1]
+ saout_R_m2_3v256x8m81_3/pcb saout_R_m2_3v256x8m81_3/vss_uq6 saout_m2_3v256x8m81_3/vdd_uq2
+ saout_R_m2_3v256x8m81_3/vdd_uq2 saout_R_m2_3v256x8m81_3/vdd_uq4 saout_R_m2_3v256x8m81_3/vdd_uq6
+ saout_R_m2_3v256x8m81_3/pcb_uq0 saout_R_m2_3v256x8m81_3/datain_uq0 saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_R_m2_3v256x8m81_3/bb[5] saout_R_m2_3v256x8m81_3/sa_3v256x8m81_0/pcb pcb[6]
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b GWE saout_R_m2_3v256x8m81_3/bb[2]
+ WEN[6] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb saout_R_m2_3v256x8m81_3/b[3]
+ saout_m2_3v256x8m81_3/ypass[7] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass saout_R_m2_3v256x8m81_3/b[6]
+ saout_R_m2_3v256x8m81_3/bb[4] saout_R_m2_3v256x8m81_3/vdd saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass
+ saout_m2_3v256x8m81_3/din_3v256x8m81_0/men saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/b
+ saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/b saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass
+ saout_R_m2_3v256x8m81_3/bb[7] saout_R_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ saout_m2_3v256x8m81_3/vdd saout_m2_3v256x8m81_3/vdd_uq0 saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass
+ VSS saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass saout_m2_3v256x8m81_3/VDD
+ saout_m2_3v256x8m81_3/vdd_uq3 saout_m2_3v256x8m81_3/VDD_uq0 saout_R_m2_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[0] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[1] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[2] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[3] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[4] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[5] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[6] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[7] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[8] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[9] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[10] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[11] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[12] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[13] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[14] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[15] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[16] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[17] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[18] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[19] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[20] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[21] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[22] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[23] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[24] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[25] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[26] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[27] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[28] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[29] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[30] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[31] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[32] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[33] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[34] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xdcap_103_novia_3v256x8m81_0[35] saout_R_m2_3v256x8m81_3/b[7] VSS saout_R_m2_3v256x8m81_3/b[7]
+ dcap_103_novia_3v256x8m81
Xsaout_m2_3v256x8m81_2 saout_m2_3v256x8m81_2/ypass[2] saout_m2_3v256x8m81_2/ypass[3]
+ saout_m2_3v256x8m81_2/ypass[4] saout_m2_3v256x8m81_2/ypass[5] saout_m2_3v256x8m81_2/ypass[6]
+ saout_m2_3v256x8m81_3/GWEN GWE saout_m2_3v256x8m81_2/bb[1] saout_m2_3v256x8m81_2/bb[4]
+ saout_m2_3v256x8m81_2/bb[7] saout_m2_3v256x8m81_2/bb[6] saout_m2_3v256x8m81_2/b[5]
+ saout_m2_3v256x8m81_2/b[7] saout_m2_3v256x8m81_2/b[2] saout_m2_3v256x8m81_2/datain
+ saout_m2_3v256x8m81_2/q saout_m2_3v256x8m81_2/pcb saout_m2_3v256x8m81_2/vss_uq4
+ saout_m2_3v256x8m81_3/vdd saout_m2_3v256x8m81_3/vdd_uq0 saout_m2_3v256x8m81_2/vdd_uq1
+ saout_m2_3v256x8m81_3/vdd_uq2 saout_m2_3v256x8m81_2/pcb_uq0 saout_m2_3v256x8m81_2/pcb_uq1
+ saout_m2_3v256x8m81_2/b[2]_uq0 saout_m2_3v256x8m81_2/b[7]_uq0 saout_m2_3v256x8m81_2/b[5]_uq0
+ saout_m2_3v256x8m81_2/bb[6]_uq0 saout_m2_3v256x8m81_2/bb[7]_uq0 saout_m2_3v256x8m81_2/bb[5]
+ saout_m2_3v256x8m81_2/bb[4]_uq0 saout_m2_3v256x8m81_2/bb[1]_uq0 saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_2/b[6] saout_m2_3v256x8m81_2/bb[2] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass
+ WEN[5] saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb saout_m2_3v256x8m81_2/b[4]
+ saout_m2_3v256x8m81_3/din_3v256x8m81_0/men GWE saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_m2_3v256x8m81_2/b[1] saout_m2_3v256x8m81_2/bb[3] saout_m2_3v256x8m81_3/ypass[7]
+ saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass
+ saout_m2_3v256x8m81_2/b[3] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass
+ saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb saout_m2_3v256x8m81_2/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ saout_m2_3v256x8m81_3/VDD_uq0 saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass
+ VSS saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ saout_m2_3v256x8m81_3/VDD saout_m2_3v256x8m81_3/vdd_uq3 saout_R_m2_3v256x8m81_3/vdd
+ saout_m2_3v256x8m81
Xsaout_m2_3v256x8m81_3 saout_m2_3v256x8m81_3/ypass[2] saout_m2_3v256x8m81_3/ypass[3]
+ saout_m2_3v256x8m81_3/ypass[4] saout_m2_3v256x8m81_3/ypass[5] saout_m2_3v256x8m81_3/ypass[6]
+ saout_m2_3v256x8m81_3/GWEN GWE saout_m2_3v256x8m81_3/bb[1] saout_m2_3v256x8m81_3/bb[4]
+ saout_m2_3v256x8m81_3/bb[7] saout_m2_3v256x8m81_3/bb[6] saout_m2_3v256x8m81_3/b[5]
+ saout_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/b[2] saout_m2_3v256x8m81_3/datain
+ saout_m2_3v256x8m81_3/q saout_m2_3v256x8m81_3/pcb saout_m2_3v256x8m81_3/vss_uq4
+ saout_m2_3v256x8m81_3/vdd saout_m2_3v256x8m81_3/vdd_uq0 saout_m2_3v256x8m81_3/vdd_uq1
+ saout_m2_3v256x8m81_3/vdd_uq2 saout_m2_3v256x8m81_3/pcb_uq0 saout_m2_3v256x8m81_3/pcb_uq1
+ saout_m2_3v256x8m81_3/b[2]_uq0 saout_m2_3v256x8m81_3/b[7]_uq0 saout_m2_3v256x8m81_3/b[5]_uq0
+ saout_m2_3v256x8m81_3/bb[6]_uq0 saout_m2_3v256x8m81_3/bb[7]_uq0 saout_m2_3v256x8m81_3/bb[5]
+ saout_m2_3v256x8m81_3/bb[4]_uq0 saout_m2_3v256x8m81_3/bb[1]_uq0 saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_3/b
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/pmos_5p0431059130201_3v256x8m81_0/D
+ saout_m2_3v256x8m81_3/b[6] saout_m2_3v256x8m81_3/bb[2] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/ypass
+ WEN[7] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/b saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/bb
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/bb saout_m2_3v256x8m81_3/b[4]
+ saout_m2_3v256x8m81_3/din_3v256x8m81_0/men GWE saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_4/b
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/ypass saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/bb
+ saout_m2_3v256x8m81_3/b[1] saout_m2_3v256x8m81_3/bb[3] saout_m2_3v256x8m81_3/ypass[7]
+ saout_R_m2_3v256x8m81_3/b[7] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_1/ypass
+ saout_m2_3v256x8m81_3/b[3] saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_5/ypass
+ saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_a_3v256x8m81_0/bb saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/bb
+ saout_m2_3v256x8m81_3/VDD_uq0 saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_2/ypass
+ VSS saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_7/ypass saout_m2_3v256x8m81_3/mux821_3v256x8m81_0/ypass_gate_3v256x8m81_6/ypass
+ saout_m2_3v256x8m81_3/VDD saout_m2_3v256x8m81_3/vdd_uq3 saout_R_m2_3v256x8m81_3/vdd
+ saout_m2_3v256x8m81
.ends

.subckt pmos_5p04310591302058_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.5499p pd=2.635u as=0.9306p ps=5.11u w=2.115u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.9306p pd=5.11u as=0.5499p ps=2.635u w=2.115u l=0.28u
.ends

.subckt pmos_1p2$$47331372_3v256x8m81 a_n42_n34# w_n133_n66# pmos_5p04310591302058_3v256x8m81_0/S_uq0
+ pmos_5p04310591302058_3v256x8m81_0/S a_118_n34# pmos_5p04310591302058_3v256x8m81_0/D
Xpmos_5p04310591302058_3v256x8m81_0 pmos_5p04310591302058_3v256x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302058_3v256x8m81_0/S_uq0 pmos_5p04310591302058_3v256x8m81_0/S
+ pmos_5p04310591302058_3v256x8m81
.ends

.subckt pmos_1p2_160_3v256x8m81 w_n133_n66# pmos_5p04310591302014_3v256x8m81_0/S pmos_5p04310591302014_3v256x8m81_0/D
+ a_n14_n34#
Xpmos_5p04310591302014_3v256x8m81_0 pmos_5p04310591302014_3v256x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302014_3v256x8m81_0/S pmos_5p04310591302014_3v256x8m81
.ends

.subckt pmos_1p2_161_3v256x8m81 pmos_5p04310591302041_3v256x8m81_0/D a_n14_89# pmos_5p04310591302041_3v256x8m81_0/S
+ w_n133_n65#
Xpmos_5p04310591302041_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_0/D a_n14_89#
+ w_n133_n65# pmos_5p04310591302041_3v256x8m81_0/S pmos_5p04310591302041_3v256x8m81
.ends

.subckt nmos_5p04310591302059_3v256x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.28u
.ends

.subckt nmos_1p2$$47329324_3v256x8m81 a_118_n34# a_n41_n34# nmos_5p04310591302059_3v256x8m81_0/S_uq0
+ nmos_5p04310591302059_3v256x8m81_0/S VSUBS nmos_5p04310591302059_3v256x8m81_0/D
Xnmos_5p04310591302059_3v256x8m81_0 nmos_5p04310591302059_3v256x8m81_0/D a_n41_n34#
+ a_118_n34# nmos_5p04310591302059_3v256x8m81_0/S_uq0 nmos_5p04310591302059_3v256x8m81_0/S
+ VSUBS nmos_5p04310591302059_3v256x8m81
.ends

.subckt nmos_1p2_157_3v256x8m81 nmos_5p04310591302010_3v256x8m81_0/D a_n14_n34# nmos_5p04310591302010_3v256x8m81_0/S
+ VSUBS
Xnmos_5p04310591302010_3v256x8m81_0 nmos_5p04310591302010_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302010_3v256x8m81_0/S VSUBS nmos_5p04310591302010_3v256x8m81
.ends

.subckt alatch_3v256x8m81 en ab a a_886_665# vdd enb vss
Xpmos_1p2$$47331372_3v256x8m81_0 nmos_5p0431059130208_3v256x8m81_1/S vdd vdd vdd nmos_5p0431059130208_3v256x8m81_1/S
+ ab pmos_1p2$$47331372_3v256x8m81
Xnmos_5p0431059130208_3v256x8m81_0 vss ab nmos_5p0431059130208_3v256x8m81_1/D vss
+ nmos_5p0431059130208_3v256x8m81
Xnmos_5p0431059130208_3v256x8m81_1 nmos_5p0431059130208_3v256x8m81_1/D enb nmos_5p0431059130208_3v256x8m81_1/S
+ vss nmos_5p0431059130208_3v256x8m81
Xpmos_1p2_160_3v256x8m81_0 vdd nmos_5p0431059130208_3v256x8m81_1/S a enb pmos_1p2_160_3v256x8m81
Xpmos_1p2_161_3v256x8m81_0 nmos_5p0431059130208_3v256x8m81_1/D a_886_665# nmos_5p0431059130208_3v256x8m81_1/S
+ vdd pmos_1p2_161_3v256x8m81
Xnmos_1p2$$47329324_3v256x8m81_0 nmos_5p0431059130208_3v256x8m81_1/S nmos_5p0431059130208_3v256x8m81_1/S
+ vss vss vss ab nmos_1p2$$47329324_3v256x8m81
Xpmos_1p2_161_3v256x8m81_1 vdd ab nmos_5p0431059130208_3v256x8m81_1/D vdd pmos_1p2_161_3v256x8m81
Xnmos_1p2_157_3v256x8m81_0 a a_886_665# nmos_5p0431059130208_3v256x8m81_1/S vss nmos_1p2_157_3v256x8m81
.ends

.subckt nmos_5p04310591302057_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.9306p pd=5.11u as=0.9306p ps=5.11u w=2.115u l=0.28u
.ends

.subckt nmos_1p2$$47514668_3v256x8m81 nmos_5p04310591302057_3v256x8m81_0/S nmos_5p04310591302057_3v256x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p04310591302057_3v256x8m81_0 nmos_5p04310591302057_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302057_3v256x8m81_0/S VSUBS nmos_5p04310591302057_3v256x8m81
.ends

.subckt ypredec1_bot_3v256x8m81 m1_n9_2295# m1_n9_2436# m1_n9_2154# alatch_3v256x8m81_0/a
+ m1_n9_2013# m1_n9_1871# pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ m1_n9_1730# pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ m3_10_2563# alatch_3v256x8m81_0/enb alatch_3v256x8m81_0/vdd VSUBS pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
Xalatch_3v256x8m81_0 alatch_3v256x8m81_0/en alatch_3v256x8m81_0/ab alatch_3v256x8m81_0/a
+ m3_10_2563# alatch_3v256x8m81_0/vdd alatch_3v256x8m81_0/enb VSUBS alatch_3v256x8m81
Xnmos_1p2$$47514668_3v256x8m81_0 VSUBS pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D VSUBS nmos_1p2$$47514668_3v256x8m81
Xnmos_1p2$$47514668_3v256x8m81_1 VSUBS pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ alatch_3v256x8m81_0/ab VSUBS nmos_1p2$$47514668_3v256x8m81
Xpmos_1p2$$46887980_3v256x8m81_0 pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D pmos_1p2$$46887980_3v256x8m81
Xpmos_1p2$$46887980_3v256x8m81_1 pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S alatch_3v256x8m81_0/ab
+ pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D pmos_1p2$$46887980_3v256x8m81
.ends

.subckt pmos_5p04310591302055_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=4.1052p pd=19.54u as=4.1052p ps=19.54u w=9.33u l=0.28u
.ends

.subckt nmos_5p04310591302054_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.8634p pd=9.35u as=1.8634p ps=9.35u w=4.235u l=0.28u
.ends

.subckt ypredec1_ys_3v256x8m81 nmos_5p04310591302054_3v256x8m81_1/D pmos_5p04310591302055_3v256x8m81_1/S
+ nmos_5p04310591302054_3v256x8m81_2/S nmos_5p04310591302054_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81_3/S
+ a_187_1127# pmos_5p04310591302055_3v256x8m81_3/D VSUBS
Xpmos_5p04310591302055_3v256x8m81_0 pmos_5p04310591302055_3v256x8m81_0/D a_187_1127#
+ pmos_5p04310591302055_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81
Xpmos_5p04310591302055_3v256x8m81_1 pmos_5p04310591302055_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81_0/D
+ pmos_5p04310591302055_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81_1/S pmos_5p04310591302055_3v256x8m81
Xpmos_5p04310591302055_3v256x8m81_2 pmos_5p04310591302055_3v256x8m81_3/S pmos_5p04310591302055_3v256x8m81_0/D
+ pmos_5p04310591302055_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81
Xpmos_5p04310591302055_3v256x8m81_3 pmos_5p04310591302055_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81_0/D
+ pmos_5p04310591302055_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81_3/S pmos_5p04310591302055_3v256x8m81
Xnmos_5p04310591302054_3v256x8m81_0 pmos_5p04310591302055_3v256x8m81_3/S pmos_5p04310591302055_3v256x8m81_0/D
+ nmos_5p04310591302054_3v256x8m81_1/D VSUBS nmos_5p04310591302054_3v256x8m81
Xnmos_5p04310591302054_3v256x8m81_1 nmos_5p04310591302054_3v256x8m81_1/D pmos_5p04310591302055_3v256x8m81_0/D
+ pmos_5p04310591302055_3v256x8m81_1/S VSUBS nmos_5p04310591302054_3v256x8m81
Xnmos_5p04310591302054_3v256x8m81_2 pmos_5p04310591302055_3v256x8m81_0/D a_187_1127#
+ nmos_5p04310591302054_3v256x8m81_2/S VSUBS nmos_5p04310591302054_3v256x8m81
Xnmos_5p04310591302054_3v256x8m81_3 nmos_5p04310591302054_3v256x8m81_3/D pmos_5p04310591302055_3v256x8m81_0/D
+ pmos_5p04310591302055_3v256x8m81_3/S VSUBS nmos_5p04310591302054_3v256x8m81
.ends

.subckt nmos_5p04310591302056_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.3916p pd=2.66u as=0.3916p ps=2.66u w=0.89u l=0.28u
.ends

.subckt nmos_5p04310591302053_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.2772p pd=2.14u as=0.2772p ps=2.14u w=0.63u l=0.28u
.ends

.subckt nmos_1p2$$47342636_3v256x8m81 nmos_5p04310591302053_3v256x8m81_0/D a_n14_n34#
+ VSUBS nmos_5p04310591302053_3v256x8m81_0/S
Xnmos_5p04310591302053_3v256x8m81_0 nmos_5p04310591302053_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302053_3v256x8m81_0/S VSUBS nmos_5p04310591302053_3v256x8m81
.ends

.subckt pmos_5p04310591302061_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=1.1836p pd=6.26u as=1.1836p ps=6.26u w=2.69u l=0.28u
.ends

.subckt pmos_1p2$$47820844_3v256x8m81 pmos_5p04310591302061_3v256x8m81_0/S a_n14_n34#
+ pmos_5p04310591302061_3v256x8m81_0/D w_n133_n65#
Xpmos_5p04310591302061_3v256x8m81_0 pmos_5p04310591302061_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302061_3v256x8m81_0/S pmos_5p04310591302061_3v256x8m81
.ends

.subckt pmos_5p04310591302060_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=1.1638p pd=6.17u as=1.1638p ps=6.17u w=2.645u l=0.28u
.ends

.subckt pmos_1p2$$47821868_3v256x8m81 pmos_5p04310591302060_3v256x8m81_0/S a_n14_n34#
+ pmos_5p04310591302060_3v256x8m81_0/D w_n133_n66#
Xpmos_5p04310591302060_3v256x8m81_0 pmos_5p04310591302060_3v256x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302060_3v256x8m81_0/S pmos_5p04310591302060_3v256x8m81
.ends

.subckt ypredec1_xa_3v256x8m81 m1_n40_n2861# a_145_n4683# m3_0_n4986# m1_n40_n3567#
+ m1_n40_n3285# pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# a_0_56# a_465_n4683# m1_n40_n3426#
+ m1_n40_n3144# pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# M3_M2$$47819820_3v256x8m81_0/VSUBS
+ pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D m1_n40_n3003#
+ a_305_n4683# pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
Xpmos_1p2$$47820844_3v256x8m81_0 pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# pmos_1p2$$47820844_3v256x8m81
Xpmos_1p2$$47820844_3v256x8m81_1 pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# pmos_1p2$$47820844_3v256x8m81
Xpmos_1p2$$47820844_3v256x8m81_2 pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# pmos_1p2$$47820844_3v256x8m81
Xpmos_1p2$$47821868_3v256x8m81_0 pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ a_145_n4683# pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D
+ pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# pmos_1p2$$47821868_3v256x8m81
Xnmos_1p2$$46551084_3v256x8m81_0 M3_M2$$47819820_3v256x8m81_0/VSUBS pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D
+ pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D M3_M2$$47819820_3v256x8m81_0/VSUBS
+ nmos_1p2$$46551084_3v256x8m81
Xnmos_1p2$$46551084_3v256x8m81_1 pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D M3_M2$$47819820_3v256x8m81_0/VSUBS
+ M3_M2$$47819820_3v256x8m81_0/VSUBS nmos_1p2$$46551084_3v256x8m81
Xpmos_1p2$$47821868_3v256x8m81_2 pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D
+ a_305_n4683# pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# pmos_1p2$$47821868_3v256x8m81
Xnmos_1p2$$46551084_3v256x8m81_2 pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D M3_M2$$47819820_3v256x8m81_0/VSUBS
+ M3_M2$$47819820_3v256x8m81_0/VSUBS nmos_1p2$$46551084_3v256x8m81
Xpmos_1p2$$47821868_3v256x8m81_3 pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ a_465_n4683# pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D
+ pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# pmos_1p2$$47821868_3v256x8m81
X0 a_361_n4624# a_305_n4683# a_201_n4624# M3_M2$$47819820_3v256x8m81_0/VSUBS nfet_03v3 ad=0.8268p pd=3.7u as=0.8268p ps=3.7u w=3.18u l=0.28u
X1 a_201_n4624# a_145_n4683# M3_M2$$47819820_3v256x8m81_0/VSUBS M3_M2$$47819820_3v256x8m81_0/VSUBS nfet_03v3 ad=0.8268p pd=3.7u as=1.4469p ps=7.27u w=3.18u l=0.28u
X2 pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/D a_465_n4683# a_361_n4624# M3_M2$$47819820_3v256x8m81_0/VSUBS nfet_03v3 ad=1.5423p pd=7.33u as=0.8268p ps=3.7u w=3.18u l=0.28u
.ends

.subckt ypredec1_xax8_3v256x8m81 ypredec1_xa_3v256x8m81_1/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_7/a_305_n4683# ypredec1_xa_3v256x8m81_6/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_2/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_7/a_465_n4683# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# ypredec1_xa_3v256x8m81_3/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# ypredec1_xa_3v256x8m81_4/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_7/a_145_n4683# ypredec1_xa_3v256x8m81_5/a_0_56# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81_5/a_465_n4683# ypredec1_xa_3v256x8m81_0/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_5/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_6/a_305_n4683# VSUBS ypredec1_xa_3v256x8m81_3/a_145_n4683#
Xypredec1_xa_3v256x8m81_0 ypredec1_xa_3v256x8m81_7/a_465_n4683# ypredec1_xa_3v256x8m81_3/a_145_n4683#
+ VSUBS ypredec1_xa_3v256x8m81_7/a_145_n4683# ypredec1_xa_3v256x8m81_5/a_465_n4683#
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# ypredec1_xa_3v256x8m81_0/a_0_56#
+ ypredec1_xa_3v256x8m81_5/a_465_n4683# ypredec1_xa_3v256x8m81_6/a_305_n4683# ypredec1_xa_3v256x8m81_3/a_145_n4683#
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# VSUBS ypredec1_xa_3v256x8m81_0/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_7/a_305_n4683# ypredec1_xa_3v256x8m81_7/a_305_n4683# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81
Xypredec1_xa_3v256x8m81_1 ypredec1_xa_3v256x8m81_7/a_465_n4683# ypredec1_xa_3v256x8m81_3/a_145_n4683#
+ VSUBS ypredec1_xa_3v256x8m81_7/a_145_n4683# ypredec1_xa_3v256x8m81_5/a_465_n4683#
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# ypredec1_xa_3v256x8m81_5/a_0_56#
+ ypredec1_xa_3v256x8m81_5/a_465_n4683# ypredec1_xa_3v256x8m81_6/a_305_n4683# ypredec1_xa_3v256x8m81_3/a_145_n4683#
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# VSUBS ypredec1_xa_3v256x8m81_1/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_7/a_305_n4683# ypredec1_xa_3v256x8m81_6/a_305_n4683# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81
Xypredec1_xa_3v256x8m81_2 ypredec1_xa_3v256x8m81_7/a_465_n4683# ypredec1_xa_3v256x8m81_3/a_145_n4683#
+ VSUBS ypredec1_xa_3v256x8m81_7/a_145_n4683# ypredec1_xa_3v256x8m81_5/a_465_n4683#
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# VSUBS ypredec1_xa_3v256x8m81_7/a_465_n4683#
+ ypredec1_xa_3v256x8m81_6/a_305_n4683# ypredec1_xa_3v256x8m81_3/a_145_n4683# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66#
+ VSUBS ypredec1_xa_3v256x8m81_2/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_7/a_305_n4683# ypredec1_xa_3v256x8m81_6/a_305_n4683# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81
Xypredec1_xa_3v256x8m81_3 ypredec1_xa_3v256x8m81_7/a_465_n4683# ypredec1_xa_3v256x8m81_3/a_145_n4683#
+ VSUBS ypredec1_xa_3v256x8m81_7/a_145_n4683# ypredec1_xa_3v256x8m81_5/a_465_n4683#
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# ypredec1_xa_3v256x8m81_3/a_0_56#
+ ypredec1_xa_3v256x8m81_7/a_465_n4683# ypredec1_xa_3v256x8m81_6/a_305_n4683# ypredec1_xa_3v256x8m81_3/a_145_n4683#
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# VSUBS ypredec1_xa_3v256x8m81_3/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_7/a_305_n4683# ypredec1_xa_3v256x8m81_7/a_305_n4683# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81
Xypredec1_xa_3v256x8m81_4 ypredec1_xa_3v256x8m81_7/a_465_n4683# ypredec1_xa_3v256x8m81_7/a_145_n4683#
+ VSUBS ypredec1_xa_3v256x8m81_7/a_145_n4683# ypredec1_xa_3v256x8m81_5/a_465_n4683#
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# ypredec1_xa_3v256x8m81_4/a_0_56#
+ ypredec1_xa_3v256x8m81_5/a_465_n4683# ypredec1_xa_3v256x8m81_6/a_305_n4683# ypredec1_xa_3v256x8m81_3/a_145_n4683#
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# VSUBS ypredec1_xa_3v256x8m81_4/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_7/a_305_n4683# ypredec1_xa_3v256x8m81_7/a_305_n4683# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81
Xypredec1_xa_3v256x8m81_5 ypredec1_xa_3v256x8m81_7/a_465_n4683# ypredec1_xa_3v256x8m81_7/a_145_n4683#
+ VSUBS ypredec1_xa_3v256x8m81_7/a_145_n4683# ypredec1_xa_3v256x8m81_5/a_465_n4683#
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# ypredec1_xa_3v256x8m81_5/a_0_56#
+ ypredec1_xa_3v256x8m81_5/a_465_n4683# ypredec1_xa_3v256x8m81_6/a_305_n4683# ypredec1_xa_3v256x8m81_3/a_145_n4683#
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# VSUBS ypredec1_xa_3v256x8m81_5/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_7/a_305_n4683# ypredec1_xa_3v256x8m81_6/a_305_n4683# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81
Xypredec1_xa_3v256x8m81_6 ypredec1_xa_3v256x8m81_7/a_465_n4683# ypredec1_xa_3v256x8m81_7/a_145_n4683#
+ VSUBS ypredec1_xa_3v256x8m81_7/a_145_n4683# ypredec1_xa_3v256x8m81_5/a_465_n4683#
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# ypredec1_xa_3v256x8m81_6/a_0_56#
+ ypredec1_xa_3v256x8m81_7/a_465_n4683# ypredec1_xa_3v256x8m81_6/a_305_n4683# ypredec1_xa_3v256x8m81_3/a_145_n4683#
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# VSUBS ypredec1_xa_3v256x8m81_6/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_7/a_305_n4683# ypredec1_xa_3v256x8m81_6/a_305_n4683# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81
Xypredec1_xa_3v256x8m81_7 ypredec1_xa_3v256x8m81_7/a_465_n4683# ypredec1_xa_3v256x8m81_7/a_145_n4683#
+ VSUBS ypredec1_xa_3v256x8m81_7/a_145_n4683# ypredec1_xa_3v256x8m81_5/a_465_n4683#
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/w_n133_n65# ypredec1_xa_3v256x8m81_7/a_0_56#
+ ypredec1_xa_3v256x8m81_7/a_465_n4683# ypredec1_xa_3v256x8m81_6/a_305_n4683# ypredec1_xa_3v256x8m81_3/a_145_n4683#
+ ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/w_n133_n66# VSUBS ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xa_3v256x8m81_7/a_305_n4683# ypredec1_xa_3v256x8m81_7/a_305_n4683# ypredec1_xa_3v256x8m81_7/pmos_1p2$$47821868_3v256x8m81_3/pmos_5p04310591302060_3v256x8m81_0/S
+ ypredec1_xa_3v256x8m81
.ends

.subckt pmos_5p04310591302062_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.2067p pd=1.315u as=0.3498p ps=2.47u w=0.795u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.3498p pd=2.47u as=0.2067p ps=1.315u w=0.795u l=0.28u
.ends

.subckt pmos_1p2$$47109164_3v256x8m81 pmos_5p04310591302062_3v256x8m81_0/S_uq0 pmos_5p04310591302062_3v256x8m81_0/D
+ pmos_5p04310591302062_3v256x8m81_0/w_n202_n86# a_118_159# pmos_5p04310591302062_3v256x8m81_0/S
+ a_n42_159#
Xpmos_5p04310591302062_3v256x8m81_0 pmos_5p04310591302062_3v256x8m81_0/D a_n42_159#
+ a_118_159# pmos_5p04310591302062_3v256x8m81_0/w_n202_n86# pmos_5p04310591302062_3v256x8m81_0/S_uq0
+ pmos_5p04310591302062_3v256x8m81_0/S pmos_5p04310591302062_3v256x8m81
.ends

.subckt ypredec1_3v256x8m81 ly[5] ly[4] ly[7] ly[2] ly[1] ly[0] ry[0] ry[1] ry[2]
+ ry[3] ry[4] ry[5] ry[6] ry[7] ly[6] men A[0] A[1] A[2] clk ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/a
+ ly[3] ypredec1_bot_3v256x8m81_0/alatch_3v256x8m81_0/a pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/w_n202_n86#
+ ypredec1_bot_3v256x8m81_1/alatch_3v256x8m81_0/a pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
Xypredec1_bot_3v256x8m81_1 ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_1/alatch_3v256x8m81_0/a ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ nmos_5p04310591302056_3v256x8m81_1/D ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb
+ ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ ypredec1_bot_3v256x8m81
Xypredec1_ys_3v256x8m81_4 M1_NWELL13_3v256x8m81_0/VSUBS ly[0] M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS ly[0] ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_5/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_bot_3v256x8m81_2 ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/a ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ nmos_5p04310591302056_3v256x8m81_1/D ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb
+ ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ ypredec1_bot_3v256x8m81
Xypredec1_ys_3v256x8m81_5 M1_NWELL13_3v256x8m81_0/VSUBS ly[1] M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS ly[1] ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_1/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_6 M1_NWELL13_3v256x8m81_0/VSUBS ly[2] M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS ly[2] ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_4/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_7 M1_NWELL13_3v256x8m81_0/VSUBS ry[5] M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS ry[5] ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_2/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_8 M1_NWELL13_3v256x8m81_0/VSUBS ry[6] M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS ry[6] ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_9 M1_NWELL13_3v256x8m81_0/VSUBS ry[7] M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS ry[7] ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_3/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_10 M1_NWELL13_3v256x8m81_0/VSUBS ry[1] M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS ry[1] ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_1/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_11 M1_NWELL13_3v256x8m81_0/VSUBS ry[2] M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS ry[2] ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_4/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_12 M1_NWELL13_3v256x8m81_0/VSUBS ry[3] M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS ry[3] ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_0/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_13 M1_NWELL13_3v256x8m81_0/VSUBS ry[4] M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS ry[4] ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_6/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xnmos_5p04310591302056_3v256x8m81_0 M1_NWELL13_3v256x8m81_0/VSUBS clk nmos_5p04310591302056_3v256x8m81_1/D
+ M1_NWELL13_3v256x8m81_0/VSUBS nmos_5p04310591302056_3v256x8m81
Xypredec1_ys_3v256x8m81_14 M1_NWELL13_3v256x8m81_0/VSUBS ry[0] M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS ry[0] ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_5/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xnmos_5p04310591302056_3v256x8m81_1 nmos_5p04310591302056_3v256x8m81_1/D men M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS nmos_5p04310591302056_3v256x8m81
Xypredec1_ys_3v256x8m81_15 M1_NWELL13_3v256x8m81_0/VSUBS ly[7] M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS ly[7] ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_3/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xnmos_1p2$$47342636_3v256x8m81_0 M1_NWELL13_3v256x8m81_0/VSUBS nmos_5p04310591302056_3v256x8m81_1/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb
+ nmos_1p2$$47342636_3v256x8m81
Xypredec1_xax8_3v256x8m81_0 ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_1/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_6/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_2/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_3/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_4/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_0/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_5/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ M1_NWELL13_3v256x8m81_0/VSUBS ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_xax8_3v256x8m81
Xypredec1_ys_3v256x8m81_0 M1_NWELL13_3v256x8m81_0/VSUBS ly[3] M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS ly[3] ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_0/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_1 M1_NWELL13_3v256x8m81_0/VSUBS ly[4] M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS ly[4] ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_6/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xypredec1_ys_3v256x8m81_2 M1_NWELL13_3v256x8m81_0/VSUBS ly[5] M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS ly[5] ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_2/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
Xpmos_1p2$$47109164_3v256x8m81_0 pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S
+ ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/w_n202_n86#
+ nmos_5p04310591302056_3v256x8m81_1/D pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S
+ nmos_5p04310591302056_3v256x8m81_1/D pmos_1p2$$47109164_3v256x8m81
Xypredec1_bot_3v256x8m81_0 ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/alatch_3v256x8m81_0/a ypredec1_bot_3v256x8m81_1/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_0/pmos_5p0431059130204_3v256x8m81_0/D
+ ypredec1_bot_3v256x8m81_0/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/D
+ nmos_5p04310591302056_3v256x8m81_1/D ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb
+ ypredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_bot_3v256x8m81_2/pmos_1p2$$46887980_3v256x8m81_1/pmos_5p0431059130204_3v256x8m81_0/S
+ ypredec1_bot_3v256x8m81
Xypredec1_ys_3v256x8m81_3 M1_NWELL13_3v256x8m81_0/VSUBS ly[6] M1_NWELL13_3v256x8m81_0/VSUBS
+ M1_NWELL13_3v256x8m81_0/VSUBS ly[6] ypredec1_xax8_3v256x8m81_0/ypredec1_xa_3v256x8m81_7/pmos_1p2$$47820844_3v256x8m81_2/pmos_5p04310591302061_3v256x8m81_0/D
+ ypredec1_ys_3v256x8m81_9/pmos_5p04310591302055_3v256x8m81_3/D M1_NWELL13_3v256x8m81_0/VSUBS
+ ypredec1_ys_3v256x8m81
X0 a_5490_186# clk nmos_5p04310591302056_3v256x8m81_1/D pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S pfet_03v3 ad=0.1917p pd=1.425u as=0.34345p ps=1.71u w=1.065u l=0.28u
X1 nmos_5p04310591302056_3v256x8m81_1/D clk a_5176_186# pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S pfet_03v3 ad=0.34345p pd=1.71u as=0.19435p ps=1.43u w=1.065u l=0.28u
X2 a_5176_186# men pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S pfet_03v3 ad=0.19435p pd=1.43u as=0.59108p ps=3.24u w=1.065u l=0.28u
X3 pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S men a_5490_186# pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/S pfet_03v3 ad=0.59108p pd=3.24u as=0.1917p ps=1.425u w=1.065u l=0.28u
.ends

.subckt pmos_5p04310591302068_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.3276p pd=11.46u as=2.3276p ps=11.46u w=5.29u l=0.28u
.ends

.subckt pmos_1p2$$47513644_3v256x8m81 pmos_5p04310591302068_3v256x8m81_0/S a_n14_n34#
+ pmos_5p04310591302068_3v256x8m81_0/D w_n133_n65#
Xpmos_5p04310591302068_3v256x8m81_0 pmos_5p04310591302068_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302068_3v256x8m81_0/S pmos_5p04310591302068_3v256x8m81
.ends

.subckt pmos_5p04310591302072_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.1406p pd=10.61u as=2.1406p ps=10.61u w=4.865u l=0.28u
.ends

.subckt pmos_1p2$$47512620_3v256x8m81 a_n14_n34# pmos_5p04310591302072_3v256x8m81_0/S
+ w_n133_n66# pmos_5p04310591302072_3v256x8m81_0/D
Xpmos_5p04310591302072_3v256x8m81_0 pmos_5p04310591302072_3v256x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302072_3v256x8m81_0/S pmos_5p04310591302072_3v256x8m81
.ends

.subckt xpredec1_xa_3v256x8m81 m1_n40_n4147# m1_n40_n4005# m3_n46_n5510# a_145_n5643#
+ m1_n40_n3864# m1_n40_n3582# m1_n40_n3723# a_0_56# m1_n40_n3441# a_465_n5643# pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/D
+ M3_M2$$47333420_3v256x8m81_1/VSUBS pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S
+ a_305_n5643#
Xpmos_1p2$$47513644_3v256x8m81_0 pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81
Xpmos_1p2$$47513644_3v256x8m81_1 pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81
Xpmos_1p2$$47513644_3v256x8m81_2 pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81
Xnmos_1p2$$47514668_3v256x8m81_0 M3_M2$$47333420_3v256x8m81_1/VSUBS pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S M3_M2$$47333420_3v256x8m81_1/VSUBS
+ nmos_1p2$$47514668_3v256x8m81
Xnmos_1p2$$47514668_3v256x8m81_1 pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/D
+ M3_M2$$47333420_3v256x8m81_1/VSUBS pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S
+ M3_M2$$47333420_3v256x8m81_1/VSUBS nmos_1p2$$47514668_3v256x8m81
Xnmos_1p2$$47514668_3v256x8m81_2 M3_M2$$47333420_3v256x8m81_1/VSUBS pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S M3_M2$$47333420_3v256x8m81_1/VSUBS
+ nmos_1p2$$47514668_3v256x8m81
Xpmos_1p2$$47512620_3v256x8m81_0 a_145_n5643# pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S
+ pmos_1p2$$47512620_3v256x8m81
Xpmos_1p2$$47512620_3v256x8m81_1 a_465_n5643# pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S
+ pmos_1p2$$47512620_3v256x8m81
Xpmos_1p2$$47512620_3v256x8m81_3 a_305_n5643# pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S
+ pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_2/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47512620_3v256x8m81
X0 a_361_n5592# a_305_n5643# a_201_n5592# M3_M2$$47333420_3v256x8m81_1/VSUBS nfet_03v3 ad=1.5145p pd=6.345u as=1.5145p ps=6.345u w=5.825u l=0.28u
X1 a_201_n5592# a_145_n5643# M3_M2$$47333420_3v256x8m81_1/VSUBS M3_M2$$47333420_3v256x8m81_1/VSUBS nfet_03v3 ad=1.5145p pd=6.345u as=2.65037p ps=12.56u w=5.825u l=0.28u
X2 pmos_1p2$$47512620_3v256x8m81_3/pmos_5p04310591302072_3v256x8m81_0/S a_465_n5643# a_361_n5592# M3_M2$$47333420_3v256x8m81_1/VSUBS nfet_03v3 ad=2.82512p pd=12.62u as=1.5145p ps=6.345u w=5.825u l=0.28u
.ends

.subckt nmos_5p04310591302071_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.3508p pd=7.02u as=1.3508p ps=7.02u w=3.07u l=0.28u
.ends

.subckt nmos_1p2$$47336492_3v256x8m81 nmos_5p04310591302071_3v256x8m81_0/S nmos_5p04310591302071_3v256x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p04310591302071_3v256x8m81_0 nmos_5p04310591302071_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302071_3v256x8m81_0/S VSUBS nmos_5p04310591302071_3v256x8m81
.ends

.subckt pmos_5p04310591302070_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=3.3528p pd=16.12u as=3.3528p ps=16.12u w=7.62u l=0.28u
.ends

.subckt pmos_1p2$$47337516_3v256x8m81 pmos_5p04310591302070_3v256x8m81_0/S pmos_5p04310591302070_3v256x8m81_0/D
+ a_n14_n34# w_n133_n65#
Xpmos_5p04310591302070_3v256x8m81_0 pmos_5p04310591302070_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302070_3v256x8m81_0/S pmos_5p04310591302070_3v256x8m81
.ends

.subckt xpredec1_bot_3v256x8m81 m1_n74_2740# pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ alatch_3v256x8m81_0/a m1_n74_3446# alatch_3v256x8m81_0/enb m1_n74_3164# m1_n74_3305#
+ m1_n74_3023# alatch_3v256x8m81_0/vdd pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/S
+ VSUBS m3_9_2964# m1_n74_2881# pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
Xnmos_1p2$$47336492_3v256x8m81_0 VSUBS pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D VSUBS nmos_1p2$$47336492_3v256x8m81
Xnmos_1p2$$47336492_3v256x8m81_1 VSUBS pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ alatch_3v256x8m81_0/ab VSUBS nmos_1p2$$47336492_3v256x8m81
Xalatch_3v256x8m81_0 alatch_3v256x8m81_0/en alatch_3v256x8m81_0/ab alatch_3v256x8m81_0/a
+ m3_9_2964# alatch_3v256x8m81_0/vdd alatch_3v256x8m81_0/enb VSUBS alatch_3v256x8m81
Xpmos_1p2$$47337516_3v256x8m81_0 pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/S
+ pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/S pmos_1p2$$47337516_3v256x8m81
Xpmos_1p2$$47337516_3v256x8m81_1 pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/S
+ pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D alatch_3v256x8m81_0/ab
+ pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/S pmos_1p2$$47337516_3v256x8m81
.ends

.subckt xpredec1_3v256x8m81 A[2] men x[7] x[6] x[5] x[4] x[3] x[2] x[1] x[0] A[1]
+ A[0] clk w_5024_6624# xpredec1_xa_3v256x8m81_7/m3_n46_n5510# pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/w_n202_n86#
+ xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd vss vdd vdd_uq0
Xxpredec1_xa_3v256x8m81_0 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/m3_n46_n5510# xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_0/a_0_56# xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ x[3] vss vdd_uq0 xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81
Xxpredec1_xa_3v256x8m81_1 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/m3_n46_n5510# xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ vss xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ x[1] vss vdd_uq0 xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81
Xxpredec1_xa_3v256x8m81_2 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/m3_n46_n5510# xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ vss xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ x[5] vss vdd_uq0 xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81
Xxpredec1_xa_3v256x8m81_3 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/m3_n46_n5510# xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_3/a_0_56# xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ x[7] vss vdd_uq0 xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81
Xxpredec1_bot_3v256x8m81_0 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ A[0] xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd vdd_uq0 vss nmos_5p04310591302056_3v256x8m81_1/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81
Xxpredec1_xa_3v256x8m81_4 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/m3_n46_n5510# xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_4/a_0_56# xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ x[2] vss vdd_uq0 xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81
Xxpredec1_bot_3v256x8m81_1 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ A[2] xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd vdd_uq0 vss nmos_5p04310591302056_3v256x8m81_1/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81
Xxpredec1_xa_3v256x8m81_5 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/m3_n46_n5510# xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_5/a_0_56# xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ x[0] vss vdd_uq0 xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81
Xxpredec1_bot_3v256x8m81_2 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ A[1] xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd vdd_uq0 vss nmos_5p04310591302056_3v256x8m81_1/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81
Xnmos_5p04310591302056_3v256x8m81_0 vss clk nmos_5p04310591302056_3v256x8m81_1/D vss
+ nmos_5p04310591302056_3v256x8m81
Xxpredec1_xa_3v256x8m81_6 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/m3_n46_n5510# xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_6/a_0_56# xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ x[4] vss vdd_uq0 xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81
Xnmos_5p04310591302056_3v256x8m81_1 nmos_5p04310591302056_3v256x8m81_1/D men vss vss
+ nmos_5p04310591302056_3v256x8m81
Xxpredec1_xa_3v256x8m81_7 xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/m3_n46_n5510# xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_0/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_0/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81_7/a_0_56# xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_bot_3v256x8m81_1/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ x[6] vss vdd_uq0 xpredec1_bot_3v256x8m81_2/pmos_1p2$$47337516_3v256x8m81_1/pmos_5p04310591302070_3v256x8m81_0/D
+ xpredec1_xa_3v256x8m81
Xnmos_1p2$$47342636_3v256x8m81_0 vss nmos_5p04310591302056_3v256x8m81_1/D vss xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb
+ nmos_1p2$$47342636_3v256x8m81
Xpmos_1p2$$47109164_3v256x8m81_0 vdd xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/enb
+ pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/w_n202_n86# nmos_5p04310591302056_3v256x8m81_1/D
+ vdd nmos_5p04310591302056_3v256x8m81_1/D pmos_1p2$$47109164_3v256x8m81
X0 a_5287_6723# men vdd w_5024_6624# pfet_03v3 ad=0.212p pd=1.46u as=0.5936p ps=3.24u w=1.06u l=0.28u
X1 a_5600_6723# clk nmos_5p04310591302056_3v256x8m81_1/D w_5024_6624# pfet_03v3 ad=0.19345p pd=1.425u as=0.32065p ps=1.665u w=1.06u l=0.28u
X2 nmos_5p04310591302056_3v256x8m81_1/D clk a_5287_6723# w_5024_6624# pfet_03v3 ad=0.32065p pd=1.665u as=0.212p ps=1.46u w=1.06u l=0.28u
X3 vdd men a_5600_6723# w_5024_6624# pfet_03v3 ad=0.5883p pd=3.23u as=0.19345p ps=1.425u w=1.06u l=0.28u
.ends

.subckt pmos_5p04310591302067_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=3.1196p pd=15.06u as=3.1196p ps=15.06u w=7.09u l=0.28u
.ends

.subckt pmos_1p2$$47643692_3v256x8m81 w_n133_n66# pmos_5p04310591302067_3v256x8m81_0/S
+ pmos_5p04310591302067_3v256x8m81_0/D a_n14_n34#
Xpmos_5p04310591302067_3v256x8m81_0 pmos_5p04310591302067_3v256x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302067_3v256x8m81_0/S pmos_5p04310591302067_3v256x8m81
.ends

.subckt nmos_1p2$$47641644_3v256x8m81 nmos_5p04310591302057_3v256x8m81_0/S nmos_5p04310591302057_3v256x8m81_0/D
+ a_n14_n34# VSUBS
Xnmos_5p04310591302057_3v256x8m81_0 nmos_5p04310591302057_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302057_3v256x8m81_0/S VSUBS nmos_5p04310591302057_3v256x8m81
.ends

.subckt pmos_1p2$$47642668_3v256x8m81 pmos_5p04310591302067_3v256x8m81_0/S pmos_5p04310591302067_3v256x8m81_0/D
+ a_n14_n34# w_n194_n66#
Xpmos_5p04310591302067_3v256x8m81_0 pmos_5p04310591302067_3v256x8m81_0/D a_n14_n34#
+ w_n194_n66# pmos_5p04310591302067_3v256x8m81_0/S pmos_5p04310591302067_3v256x8m81
.ends

.subckt xpredec0_xa_3v256x8m81 m3_107_5938# m1_255_3759# a_612_1974# m1_255_3263#
+ m1_255_3619# m1_255_3901# m3_598_2319# pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D
+ a_472_3898# M3_M2$$47644716_3v256x8m81_2/VSUBS pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D
+ nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S nmos_1p2$$47641644_3v256x8m81_3/nmos_5p04310591302057_3v256x8m81_0/D
+ pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/S
Xpmos_1p2$$47513644_3v256x8m81_0 pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D pmos_1p2$$47513644_3v256x8m81
Xpmos_1p2$$47513644_3v256x8m81_1 pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D pmos_1p2$$47513644_3v256x8m81
Xpmos_1p2$$47513644_3v256x8m81_2 pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D pmos_1p2$$47513644_3v256x8m81
Xpmos_1p2$$47513644_3v256x8m81_3 pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/S
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D pmos_1p2$$47513644_3v256x8m81
Xpmos_1p2$$47643692_3v256x8m81_0 pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D
+ a_472_3898# pmos_1p2$$47643692_3v256x8m81
Xnmos_1p2$$47641644_3v256x8m81_0 nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S
+ M3_M2$$47644716_3v256x8m81_2/VSUBS nmos_1p2$$47641644_3v256x8m81
Xnmos_1p2$$47641644_3v256x8m81_1 nmos_1p2$$47641644_3v256x8m81_3/nmos_5p04310591302057_3v256x8m81_0/D
+ pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S
+ M3_M2$$47644716_3v256x8m81_2/VSUBS nmos_1p2$$47641644_3v256x8m81
Xpmos_1p2$$47642668_3v256x8m81_0 pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S a_612_1974#
+ pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/D pmos_1p2$$47642668_3v256x8m81
Xnmos_1p2$$47641644_3v256x8m81_2 pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D
+ nmos_1p2$$47641644_3v256x8m81_3/nmos_5p04310591302057_3v256x8m81_0/D pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S
+ M3_M2$$47644716_3v256x8m81_2/VSUBS nmos_1p2$$47641644_3v256x8m81
Xnmos_1p2$$47641644_3v256x8m81_3 pmos_1p2$$47513644_3v256x8m81_3/pmos_5p04310591302068_3v256x8m81_0/D
+ nmos_1p2$$47641644_3v256x8m81_3/nmos_5p04310591302057_3v256x8m81_0/D pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S
+ M3_M2$$47644716_3v256x8m81_2/VSUBS nmos_1p2$$47641644_3v256x8m81
X0 M3_M2$$47644716_3v256x8m81_2/VSUBS a_612_1974# a_539_2025# M3_M2$$47644716_3v256x8m81_2/VSUBS nfet_03v3 ad=3.1746p pd=12.55u as=1.0439p ps=6.085u w=5.72u l=0.28u
X1 a_539_2025# a_472_3898# pmos_1p2$$47643692_3v256x8m81_0/pmos_5p04310591302067_3v256x8m81_0/S M3_M2$$47644716_3v256x8m81_2/VSUBS nfet_03v3 ad=1.0439p pd=6.085u as=3.146p ps=12.54u w=5.72u l=0.28u
.ends

.subckt pmos_5p04310591302063_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=2.7016p pd=13.16u as=2.7016p ps=13.16u w=6.14u l=0.28u
.ends

.subckt pmos_1p2$$47504428_3v256x8m81 a_n14_n34# pmos_5p04310591302063_3v256x8m81_0/D
+ w_n133_n66# pmos_5p04310591302063_3v256x8m81_0/S
Xpmos_5p04310591302063_3v256x8m81_0 pmos_5p04310591302063_3v256x8m81_0/D a_n14_n34#
+ w_n133_n66# pmos_5p04310591302063_3v256x8m81_0/S pmos_5p04310591302063_3v256x8m81
.ends

.subckt nmos_5p04310591302065_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.0714p pd=5.75u as=1.0714p ps=5.75u w=2.435u l=0.28u
.ends

.subckt nmos_1p2$$47502380_3v256x8m81 nmos_5p04310591302065_3v256x8m81_0/S a_n14_n34#
+ nmos_5p04310591302065_3v256x8m81_0/D VSUBS
Xnmos_5p04310591302065_3v256x8m81_0 nmos_5p04310591302065_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302065_3v256x8m81_0/S VSUBS nmos_5p04310591302065_3v256x8m81
.ends

.subckt pmos_5p04310591302064_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=3.6322p pd=17.39u as=3.6322p ps=17.39u w=8.255u l=0.28u
.ends

.subckt pmos_1p2$$47503404_3v256x8m81 pmos_5p04310591302064_3v256x8m81_0/S a_n14_n34#
+ pmos_5p04310591302064_3v256x8m81_0/D w_n133_n65#
Xpmos_5p04310591302064_3v256x8m81_0 pmos_5p04310591302064_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302064_3v256x8m81_0/S pmos_5p04310591302064_3v256x8m81
.ends

.subckt nmos_5p04310591302066_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.4454p pd=7.45u as=1.4454p ps=7.45u w=3.285u l=0.28u
.ends

.subckt xpredec0_bot_3v256x8m81 nmos_5p04310591302066_3v256x8m81_0/D nmos_1p2$$47502380_3v256x8m81_0/nmos_5p04310591302065_3v256x8m81_0/S
+ pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D m1_n74_3354#
+ m1_n74_3071# m1_n74_3213# alatch_3v256x8m81_0/a alatch_3v256x8m81_0/vdd m1_n74_2930#
+ VSUBS m3_10_3351# alatch_3v256x8m81_0/enb pmos_1p2$$47503404_3v256x8m81_0/pmos_5p04310591302064_3v256x8m81_0/S
+ pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/S
Xpmos_1p2$$47504428_3v256x8m81_0 nmos_5p04310591302066_3v256x8m81_0/D pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ pmos_1p2$$47503404_3v256x8m81_0/pmos_5p04310591302064_3v256x8m81_0/S pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/S
+ pmos_1p2$$47504428_3v256x8m81
Xnmos_1p2$$47502380_3v256x8m81_0 nmos_1p2$$47502380_3v256x8m81_0/nmos_5p04310591302065_3v256x8m81_0/S
+ nmos_5p04310591302066_3v256x8m81_0/D pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ VSUBS nmos_1p2$$47502380_3v256x8m81
Xalatch_3v256x8m81_0 alatch_3v256x8m81_0/en alatch_3v256x8m81_0/ab alatch_3v256x8m81_0/a
+ m3_10_3351# alatch_3v256x8m81_0/vdd alatch_3v256x8m81_0/enb VSUBS alatch_3v256x8m81
Xpmos_1p2$$47503404_3v256x8m81_0 pmos_1p2$$47503404_3v256x8m81_0/pmos_5p04310591302064_3v256x8m81_0/S
+ alatch_3v256x8m81_0/ab nmos_5p04310591302066_3v256x8m81_0/D pmos_1p2$$47503404_3v256x8m81_0/pmos_5p04310591302064_3v256x8m81_0/S
+ pmos_1p2$$47503404_3v256x8m81
Xnmos_5p04310591302066_3v256x8m81_0 nmos_5p04310591302066_3v256x8m81_0/D alatch_3v256x8m81_0/ab
+ VSUBS VSUBS nmos_5p04310591302066_3v256x8m81
.ends

.subckt pmos_5p04310591302069_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.1378p pd=1.05u as=0.2332p ps=1.94u w=0.53u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.2332p pd=1.94u as=0.1378p ps=1.05u w=0.53u l=0.28u
.ends

.subckt xpredec0_3v256x8m81 vss A[0] x[0] x[1] x[2] x[3] A[1] clk vss_uq0 vdd_uq0
+ men vdd xpredec0_xa_3v256x8m81_3/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ xpredec0_xa_3v256x8m81_2/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ VSUBS vdd_uq2
Xxpredec0_xa_3v256x8m81_3 VSUBS xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D
+ vdd vdd_uq2 xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D VSUBS
+ x[3] xpredec0_xa_3v256x8m81_3/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ VSUBS vdd_uq2 xpredec0_xa_3v256x8m81
Xnmos_5p04310591302040_3v256x8m81_0 nmos_5p04310591302040_3v256x8m81_1/S men VSUBS
+ VSUBS nmos_5p04310591302040_3v256x8m81
Xnmos_5p04310591302040_3v256x8m81_1 VSUBS clk nmos_5p04310591302040_3v256x8m81_1/S
+ VSUBS nmos_5p04310591302040_3v256x8m81
Xxpredec0_bot_3v256x8m81_0 xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D
+ VSUBS xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ A[0] vdd xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ VSUBS nmos_5p04310591302040_3v256x8m81_1/S pmos_5p04310591302069_3v256x8m81_0/D
+ vdd_uq2 vdd_uq2 xpredec0_bot_3v256x8m81
Xnmos_1p2$$46563372_3v256x8m81_0 VSUBS nmos_5p04310591302040_3v256x8m81_1/S pmos_5p04310591302069_3v256x8m81_0/D
+ VSUBS nmos_1p2$$46563372_3v256x8m81
Xxpredec0_bot_3v256x8m81_1 xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D
+ VSUBS xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ A[1] vdd xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ VSUBS nmos_5p04310591302040_3v256x8m81_1/S pmos_5p04310591302069_3v256x8m81_0/D
+ vdd_uq2 vdd_uq2 xpredec0_bot_3v256x8m81
Xxpredec0_xa_3v256x8m81_0 VSUBS xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D
+ vdd vdd_uq2 xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ VSUBS x[0] xpredec0_xa_3v256x8m81_2/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ VSUBS vdd_uq2 xpredec0_xa_3v256x8m81
Xxpredec0_xa_3v256x8m81_1 VSUBS xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D
+ vdd vdd_uq2 xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D VSUBS
+ x[2] xpredec0_xa_3v256x8m81_3/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ VSUBS vdd_uq2 xpredec0_xa_3v256x8m81
Xpmos_5p04310591302069_3v256x8m81_0 pmos_5p04310591302069_3v256x8m81_0/D nmos_5p04310591302040_3v256x8m81_1/S
+ nmos_5p04310591302040_3v256x8m81_1/S vdd_uq2 vdd_uq2 vdd_uq2 pmos_5p04310591302069_3v256x8m81
Xxpredec0_xa_3v256x8m81_2 VSUBS xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D xpredec0_bot_3v256x8m81_0/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ xpredec0_bot_3v256x8m81_0/nmos_5p04310591302066_3v256x8m81_0/D xpredec0_bot_3v256x8m81_1/nmos_5p04310591302066_3v256x8m81_0/D
+ vdd vdd_uq2 xpredec0_bot_3v256x8m81_1/pmos_1p2$$47504428_3v256x8m81_0/pmos_5p04310591302063_3v256x8m81_0/D
+ VSUBS x[1] xpredec0_xa_3v256x8m81_2/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ VSUBS vdd_uq2 xpredec0_xa_3v256x8m81
X0 vdd_uq2 men a_3416_6773# vdd_uq2 pfet_03v3 ad=0.448p pd=2.72u as=0.162p ps=1.205u w=0.8u l=0.28u
X1 nmos_5p04310591302040_3v256x8m81_1/S clk a_3091_6773# vdd_uq2 pfet_03v3 ad=0.218p pd=1.345u as=0.208p ps=1.32u w=0.8u l=0.28u
X2 a_3091_6773# men vdd_uq2 vdd_uq2 pfet_03v3 ad=0.208p pd=1.32u as=0.364p ps=2.51u w=0.8u l=0.28u
X3 a_3416_6773# clk nmos_5p04310591302040_3v256x8m81_1/S vdd_uq2 pfet_03v3 ad=0.162p pd=1.205u as=0.218p ps=1.345u w=0.8u l=0.28u
.ends

.subckt prexdec_top_3v256x8m81 A[2] A[6] xb[3] xc[1] xc[2] xc[3] xb[1] xb[2] xb[0]
+ xa[1] xa[2] xa[4] xa[5] xa[6] xa[7] A[0] A[3] A[5] A[1] xa[0] xpredec0_3v256x8m81_1/xpredec0_xa_3v256x8m81_3/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ xa[3] xpredec1_3v256x8m81_0/clk xpredec0_3v256x8m81_0/xpredec0_xa_3v256x8m81_3/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ xpredec0_3v256x8m81_1/xpredec0_xa_3v256x8m81_2/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ xpredec1_3v256x8m81_0/w_5024_6624# xpredec0_3v256x8m81_0/xpredec0_xa_3v256x8m81_2/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ xpredec1_3v256x8m81_0/pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/w_n202_n86#
+ A[4] xc[0] men xpredec0_3v256x8m81_1/vdd xpredec1_3v256x8m81_0/xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd
+ xpredec0_3v256x8m81_1/clk xpredec1_3v256x8m81_0/vdd VSUBS
Xxpredec1_3v256x8m81_0 A[2] men xa[7] xa[6] xa[5] xa[4] xa[3] xa[2] xa[1] xa[0] A[1]
+ A[0] xpredec1_3v256x8m81_0/clk xpredec1_3v256x8m81_0/w_5024_6624# xpredec0_3v256x8m81_1/vdd
+ xpredec1_3v256x8m81_0/pmos_1p2$$47109164_3v256x8m81_0/pmos_5p04310591302062_3v256x8m81_0/w_n202_n86#
+ xpredec1_3v256x8m81_0/xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd VSUBS xpredec1_3v256x8m81_0/vdd
+ xpredec1_3v256x8m81_0/vdd xpredec1_3v256x8m81
Xxpredec0_3v256x8m81_0 xpredec0_3v256x8m81_0/vss A[3] xb[0] xb[1] xb[2] xb[3] A[4]
+ xpredec0_3v256x8m81_1/clk xpredec0_3v256x8m81_0/vss_uq0 xpredec0_3v256x8m81_0/vdd_uq0
+ men xpredec0_3v256x8m81_1/vdd xpredec0_3v256x8m81_0/xpredec0_xa_3v256x8m81_3/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ xpredec0_3v256x8m81_0/xpredec0_xa_3v256x8m81_2/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ VSUBS xpredec1_3v256x8m81_0/vdd xpredec0_3v256x8m81
Xxpredec0_3v256x8m81_1 VSUBS A[5] xc[0] xc[1] xc[2] xc[3] A[6] xpredec0_3v256x8m81_1/clk
+ VSUBS xpredec0_3v256x8m81_1/vdd men xpredec0_3v256x8m81_1/vdd xpredec0_3v256x8m81_1/xpredec0_xa_3v256x8m81_3/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ xpredec0_3v256x8m81_1/xpredec0_xa_3v256x8m81_2/nmos_1p2$$47641644_3v256x8m81_0/nmos_5p04310591302057_3v256x8m81_0/S
+ VSUBS xpredec1_3v256x8m81_0/vdd xpredec0_3v256x8m81
.ends

.subckt pmos_5p04310591302088_3v256x8m81 D_uq2 D_uq1 D_uq0 D a_n252_n44# a_550_n44#
+ a_229_n44# w_n426_n86# S_uq4 S_uq2 S_uq3 S_uq1 a_390_n44# S_uq0 S a_n92_n44# a_1032_n44#
+ a_1192_n44# a_711_n44# a_69_n44# D_uq3 a_871_n44#
X0 D_uq1 a_390_n44# S_uq2 w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=1.52775p ps=6.345u w=5.82u l=0.28u
X1 D_uq3 a_n252_n44# S_uq4 w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=2.5608p ps=12.52u w=5.82u l=0.28u
X2 D_uq2 a_69_n44# S_uq3 w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=1.52775p ps=6.345u w=5.82u l=0.28u
X3 S_uq2 a_229_n44# D_uq2 w_n426_n86# pfet_03v3 ad=1.52775p pd=6.345u as=1.5132p ps=6.34u w=5.82u l=0.28u
X4 S_uq1 a_550_n44# D_uq1 w_n426_n86# pfet_03v3 ad=1.52775p pd=6.345u as=1.5132p ps=6.34u w=5.82u l=0.28u
X5 S_uq0 a_1192_n44# D_uq0 w_n426_n86# pfet_03v3 ad=2.5608p pd=12.52u as=1.5132p ps=6.34u w=5.82u l=0.28u
X6 D_uq0 a_1032_n44# S w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=1.52775p ps=6.345u w=5.82u l=0.28u
X7 S_uq3 a_n92_n44# D_uq3 w_n426_n86# pfet_03v3 ad=1.52775p pd=6.345u as=1.5132p ps=6.34u w=5.82u l=0.28u
X8 S a_871_n44# D w_n426_n86# pfet_03v3 ad=1.52775p pd=6.345u as=1.5132p ps=6.34u w=5.82u l=0.28u
X9 D a_711_n44# S_uq1 w_n426_n86# pfet_03v3 ad=1.5132p pd=6.34u as=1.52775p ps=6.345u w=5.82u l=0.28u
.ends

.subckt nmos_5p04310591302081_3v256x8m81 D_uq2 D_uq1 D_uq0 D a_634_n44# a_n168_n44#
+ a_313_n44# a_795_n44# S_uq2 a_474_n44# S_uq1 a_n8_n44# S_uq0 S a_153_n44# VSUBS
X0 D_uq1 a_153_n44# S_uq1 VSUBS nfet_03v3 ad=0.1079p pd=0.935u as=0.10892p ps=0.94u w=0.415u l=0.28u
X1 D a_474_n44# S VSUBS nfet_03v3 ad=0.1079p pd=0.935u as=0.10892p ps=0.94u w=0.415u l=0.28u
X2 D_uq2 a_n168_n44# S_uq2 VSUBS nfet_03v3 ad=0.1079p pd=0.935u as=0.1826p ps=1.71u w=0.415u l=0.28u
X3 S_uq1 a_n8_n44# D_uq2 VSUBS nfet_03v3 ad=0.10892p pd=0.94u as=0.1079p ps=0.935u w=0.415u l=0.28u
X4 D_uq0 a_795_n44# S_uq0 VSUBS nfet_03v3 ad=0.1826p pd=1.71u as=0.10892p ps=0.94u w=0.415u l=0.28u
X5 S a_313_n44# D_uq1 VSUBS nfet_03v3 ad=0.10892p pd=0.94u as=0.1079p ps=0.935u w=0.415u l=0.28u
X6 S_uq0 a_634_n44# D VSUBS nfet_03v3 ad=0.10892p pd=0.94u as=0.1079p ps=0.935u w=0.415u l=0.28u
.ends

.subckt pmos_5p04310591302077_3v256x8m81 D_uq2 D_uq1 D_uq0 D a_n252_n44# a_550_n44#
+ a_229_n44# w_n426_n86# S_uq4 S_uq2 S_uq3 S_uq1 a_390_n44# S_uq0 S a_n92_n44# a_1032_n44#
+ a_1192_n44# a_711_n44# a_69_n44# D_uq3 a_871_n44#
X0 D_uq1 a_390_n44# S_uq2 w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.5775p ps=2.725u w=2.2u l=0.28u
X1 D_uq3 a_n252_n44# S_uq4 w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.968p ps=5.28u w=2.2u l=0.28u
X2 D_uq2 a_69_n44# S_uq3 w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.5775p ps=2.725u w=2.2u l=0.28u
X3 S_uq2 a_229_n44# D_uq2 w_n426_n86# pfet_03v3 ad=0.5775p pd=2.725u as=0.572p ps=2.72u w=2.2u l=0.28u
X4 S_uq1 a_550_n44# D_uq1 w_n426_n86# pfet_03v3 ad=0.5775p pd=2.725u as=0.572p ps=2.72u w=2.2u l=0.28u
X5 S_uq0 a_1192_n44# D_uq0 w_n426_n86# pfet_03v3 ad=0.968p pd=5.28u as=0.572p ps=2.72u w=2.2u l=0.28u
X6 D_uq0 a_1032_n44# S w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.5775p ps=2.725u w=2.2u l=0.28u
X7 S_uq3 a_n92_n44# D_uq3 w_n426_n86# pfet_03v3 ad=0.5775p pd=2.725u as=0.572p ps=2.72u w=2.2u l=0.28u
X8 S a_871_n44# D w_n426_n86# pfet_03v3 ad=0.5775p pd=2.725u as=0.572p ps=2.72u w=2.2u l=0.28u
X9 D a_711_n44# S_uq1 w_n426_n86# pfet_03v3 ad=0.572p pd=2.72u as=0.5775p ps=2.725u w=2.2u l=0.28u
.ends

.subckt nmos_5p04310591302075_3v256x8m81 D_uq2 D_uq1 D_uq0 D a_n252_n44# a_550_n44#
+ a_229_n44# S_uq4 S_uq2 S_uq3 S_uq1 a_390_n44# S_uq0 S a_n92_n44# a_1032_n44# a_1192_n44#
+ a_711_n44# a_69_n44# D_uq3 a_871_n44# VSUBS
X0 D_uq1 a_390_n44# S_uq2 VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.23492p ps=1.42u w=0.895u l=0.28u
X1 D_uq3 a_n252_n44# S_uq4 VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.3938p ps=2.67u w=0.895u l=0.28u
X2 D_uq2 a_69_n44# S_uq3 VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.23492p ps=1.42u w=0.895u l=0.28u
X3 S_uq2 a_229_n44# D_uq2 VSUBS nfet_03v3 ad=0.23492p pd=1.42u as=0.2327p ps=1.415u w=0.895u l=0.28u
X4 S_uq1 a_550_n44# D_uq1 VSUBS nfet_03v3 ad=0.23492p pd=1.42u as=0.2327p ps=1.415u w=0.895u l=0.28u
X5 S_uq0 a_1192_n44# D_uq0 VSUBS nfet_03v3 ad=0.3938p pd=2.67u as=0.2327p ps=1.415u w=0.895u l=0.28u
X6 D_uq0 a_1032_n44# S VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.23492p ps=1.42u w=0.895u l=0.28u
X7 S_uq3 a_n92_n44# D_uq3 VSUBS nfet_03v3 ad=0.23492p pd=1.42u as=0.2327p ps=1.415u w=0.895u l=0.28u
X8 S a_871_n44# D VSUBS nfet_03v3 ad=0.23492p pd=1.42u as=0.2327p ps=1.415u w=0.895u l=0.28u
X9 D a_711_n44# S_uq1 VSUBS nfet_03v3 ad=0.2327p pd=1.415u as=0.23492p ps=1.42u w=0.895u l=0.28u
.ends

.subckt pmos_5p04310591302080_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.3445p pd=1.845u as=0.583p ps=3.53u w=1.325u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.583p pd=3.53u as=0.3445p ps=1.845u w=1.325u l=0.28u
.ends

.subckt nmos_5p04310591302076_3v256x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.28u
.ends

.subckt pmos_5p04310591302079_3v256x8m81 D_uq2 D_uq1 D_uq0 D a_486_n44# a_165_n44#
+ a_n156_n44# S_uq2 S_uq1 S_uq0 S a_4_n44# a_646_n44# w_n330_n86# a_808_n44# a_325_n44#
X0 S_uq0 a_646_n44# D w_n330_n86# pfet_03v3 ad=0.27162p pd=1.555u as=0.2665p ps=1.545u w=1.025u l=0.28u
X1 D_uq1 a_165_n44# S_uq1 w_n330_n86# pfet_03v3 ad=0.2665p pd=1.545u as=0.26905p ps=1.55u w=1.025u l=0.28u
X2 D a_486_n44# S w_n330_n86# pfet_03v3 ad=0.2665p pd=1.545u as=0.26905p ps=1.55u w=1.025u l=0.28u
X3 S_uq1 a_4_n44# D_uq2 w_n330_n86# pfet_03v3 ad=0.26905p pd=1.55u as=0.2665p ps=1.545u w=1.025u l=0.28u
X4 D_uq2 a_n156_n44# S_uq2 w_n330_n86# pfet_03v3 ad=0.2665p pd=1.545u as=0.451p ps=2.93u w=1.025u l=0.28u
X5 S a_325_n44# D_uq1 w_n330_n86# pfet_03v3 ad=0.26905p pd=1.55u as=0.2665p ps=1.545u w=1.025u l=0.28u
X6 D_uq0 a_808_n44# S_uq0 w_n330_n86# pfet_03v3 ad=0.451p pd=2.93u as=0.27162p ps=1.555u w=1.025u l=0.28u
.ends

.subckt pmos_5p04310591302082_3v256x8m81 a_20_n44# D_uq1 D_uq0 D a_181_n44# a_502_n44#
+ S_uq2 a_662_n44# S_uq1 a_n140_n44# S_uq0 S a_341_n44# w_n314_n86#
X0 S a_341_n44# D w_n314_n86# pfet_03v3 ad=0.30318p pd=1.68u as=0.3003p ps=1.675u w=1.155u l=0.28u
X1 S_uq0 a_662_n44# D_uq0 w_n314_n86# pfet_03v3 ad=0.5082p pd=3.19u as=0.3003p ps=1.675u w=1.155u l=0.28u
X2 D_uq0 a_502_n44# S w_n314_n86# pfet_03v3 ad=0.3003p pd=1.675u as=0.30318p ps=1.68u w=1.155u l=0.28u
X3 S_uq1 a_20_n44# D_uq1 w_n314_n86# pfet_03v3 ad=0.30318p pd=1.68u as=0.3003p ps=1.675u w=1.155u l=0.28u
X4 D a_181_n44# S_uq1 w_n314_n86# pfet_03v3 ad=0.3003p pd=1.675u as=0.30318p ps=1.68u w=1.155u l=0.28u
X5 D_uq1 a_n140_n44# S_uq2 w_n314_n86# pfet_03v3 ad=0.3003p pd=1.675u as=0.5082p ps=3.19u w=1.155u l=0.28u
.ends

.subckt nmos_5p04310591302078_3v256x8m81 D_uq0 D S_uq0 S a_217_n44# a_n104_n44# a_56_n44#
+ VSUBS
X0 D_uq0 a_217_n44# S_uq0 VSUBS nfet_03v3 ad=0.4092p pd=2.74u as=0.24412p ps=1.455u w=0.93u l=0.28u
X1 S_uq0 a_56_n44# D VSUBS nfet_03v3 ad=0.24412p pd=1.455u as=0.2418p ps=1.45u w=0.93u l=0.28u
X2 D a_n104_n44# S VSUBS nfet_03v3 ad=0.2418p pd=1.45u as=0.4092p ps=2.74u w=0.93u l=0.28u
.ends

.subckt wen_v2_3v256x8m81 clk wen GWE vdd IGWEN vss
Xnmos_1p2$$202596396_3v256x8m81_0 vss pmos_5p04310591302014_3v256x8m81_2/S pmos_5p04310591302041_3v256x8m81_1/D
+ vss nmos_1p2$$202596396_3v256x8m81
Xpmos_5p04310591302041_3v256x8m81_0 nmos_5p0431059130208_3v256x8m81_1/D nmos_5p0431059130208_3v256x8m81_4/D
+ vdd nmos_5p0431059130208_3v256x8m81_1/S pmos_5p04310591302041_3v256x8m81
Xpmos_5p04310591302041_3v256x8m81_1 pmos_5p04310591302041_3v256x8m81_1/D nmos_5p0431059130208_3v256x8m81_3/D
+ vdd pmos_5p04310591302041_3v256x8m81_1/S pmos_5p04310591302041_3v256x8m81
Xnmos_5p04310591302081_3v256x8m81_0 pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D
+ pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D nmos_5p0431059130208_3v256x8m81_1/S
+ nmos_5p0431059130208_3v256x8m81_1/S nmos_5p0431059130208_3v256x8m81_1/S nmos_5p0431059130208_3v256x8m81_1/S
+ vss nmos_5p0431059130208_3v256x8m81_1/S vss nmos_5p0431059130208_3v256x8m81_1/S
+ vss vss nmos_5p0431059130208_3v256x8m81_1/S vss nmos_5p04310591302081_3v256x8m81
Xpmos_5p04310591302077_3v256x8m81_0 IGWEN IGWEN IGWEN IGWEN pmos_5p04310591302082_3v256x8m81_0/D
+ pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D vdd vdd
+ vdd vdd vdd pmos_5p04310591302082_3v256x8m81_0/D vdd vdd pmos_5p04310591302082_3v256x8m81_0/D
+ pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D
+ pmos_5p04310591302082_3v256x8m81_0/D IGWEN pmos_5p04310591302082_3v256x8m81_0/D
+ pmos_5p04310591302077_3v256x8m81
Xpmos_5p04310591302077_3v256x8m81_2 GWE GWE GWE GWE pmos_5p04310591302079_3v256x8m81_0/D
+ pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D vdd vdd
+ vdd vdd vdd pmos_5p04310591302079_3v256x8m81_0/D vdd vdd pmos_5p04310591302079_3v256x8m81_0/D
+ pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D
+ pmos_5p04310591302079_3v256x8m81_0/D GWE pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302077_3v256x8m81
Xnmos_5p04310591302075_3v256x8m81_0 GWE GWE GWE GWE pmos_5p04310591302079_3v256x8m81_0/D
+ pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D vss vss
+ vss vss pmos_5p04310591302079_3v256x8m81_0/D vss vss pmos_5p04310591302079_3v256x8m81_0/D
+ pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D
+ pmos_5p04310591302079_3v256x8m81_0/D GWE pmos_5p04310591302079_3v256x8m81_0/D vss
+ nmos_5p04310591302075_3v256x8m81
Xnmos_5p0431059130208_3v256x8m81_0 vss pmos_5p04310591302079_3v256x8m81_0/D nmos_5p0431059130208_3v256x8m81_1/D
+ vss nmos_5p0431059130208_3v256x8m81
Xnmos_5p04310591302075_3v256x8m81_1 IGWEN IGWEN IGWEN IGWEN pmos_5p04310591302082_3v256x8m81_0/D
+ pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D vss vss
+ vss vss pmos_5p04310591302082_3v256x8m81_0/D vss vss pmos_5p04310591302082_3v256x8m81_0/D
+ pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D
+ pmos_5p04310591302082_3v256x8m81_0/D IGWEN pmos_5p04310591302082_3v256x8m81_0/D
+ vss nmos_5p04310591302075_3v256x8m81
Xnmos_5p0431059130208_3v256x8m81_1 nmos_5p0431059130208_3v256x8m81_1/D nmos_5p0431059130208_3v256x8m81_3/D
+ nmos_5p0431059130208_3v256x8m81_1/S vss nmos_5p0431059130208_3v256x8m81
Xpmos_5p04310591302080_3v256x8m81_0 pmos_5p04310591302080_3v256x8m81_0/D pmos_5p04310591302014_3v256x8m81_2/S
+ pmos_5p04310591302014_3v256x8m81_2/S vdd vdd vdd pmos_5p04310591302080_3v256x8m81
Xnmos_5p0431059130208_3v256x8m81_2 vss wen nmos_5p0431059130208_3v256x8m81_2/S vss
+ nmos_5p0431059130208_3v256x8m81
Xnmos_5p0431059130208_3v256x8m81_3 nmos_5p0431059130208_3v256x8m81_3/D clk vss vss
+ nmos_5p0431059130208_3v256x8m81
Xnmos_5p0431059130208_3v256x8m81_4 nmos_5p0431059130208_3v256x8m81_4/D nmos_5p0431059130208_3v256x8m81_3/D
+ vss vss nmos_5p0431059130208_3v256x8m81
Xnmos_5p04310591302010_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_1/S nmos_5p0431059130208_3v256x8m81_3/D
+ nmos_5p0431059130208_3v256x8m81_2/S vss nmos_5p04310591302010_3v256x8m81
Xnmos_5p04310591302076_3v256x8m81_0 pmos_5p04310591302080_3v256x8m81_0/D pmos_5p04310591302014_3v256x8m81_2/S
+ pmos_5p04310591302014_3v256x8m81_2/S vss vss vss nmos_5p04310591302076_3v256x8m81
Xpmos_1p2$$202587180_3v256x8m81_0 nmos_5p0431059130208_3v256x8m81_2/S nmos_5p0431059130208_3v256x8m81_4/D
+ pmos_5p04310591302041_3v256x8m81_1/S vdd pmos_1p2$$202587180_3v256x8m81
Xpmos_5p04310591302079_3v256x8m81_0 pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D
+ pmos_5p04310591302079_3v256x8m81_0/D pmos_5p04310591302079_3v256x8m81_0/D nmos_5p0431059130208_3v256x8m81_1/S
+ nmos_5p0431059130208_3v256x8m81_1/S nmos_5p0431059130208_3v256x8m81_1/S vdd vdd
+ vdd vdd nmos_5p0431059130208_3v256x8m81_1/S nmos_5p0431059130208_3v256x8m81_1/S
+ vdd nmos_5p0431059130208_3v256x8m81_1/S nmos_5p0431059130208_3v256x8m81_1/S pmos_5p04310591302079_3v256x8m81
Xpmos_5p04310591302020_3v256x8m81_0 pmos_5p04310591302080_3v256x8m81_0/D nmos_5p0431059130208_3v256x8m81_3/D
+ nmos_5p0431059130208_3v256x8m81_3/D vdd nmos_5p0431059130208_3v256x8m81_1/S nmos_5p0431059130208_3v256x8m81_1/S
+ pmos_5p04310591302020_3v256x8m81
Xnmos_5p04310591302039_3v256x8m81_0 pmos_5p04310591302080_3v256x8m81_0/D nmos_5p0431059130208_3v256x8m81_4/D
+ nmos_5p0431059130208_3v256x8m81_4/D nmos_5p0431059130208_3v256x8m81_1/S nmos_5p0431059130208_3v256x8m81_1/S
+ vss nmos_5p04310591302039_3v256x8m81
Xpmos_1p2$$202586156_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_1/D pmos_5p04310591302014_3v256x8m81_2/S
+ vdd vdd pmos_1p2$$202586156_3v256x8m81
Xnmos_1p2$$202595372_3v256x8m81_0 vss pmos_5p04310591302041_3v256x8m81_1/S pmos_5p04310591302014_3v256x8m81_2/S
+ vss nmos_1p2$$202595372_3v256x8m81
Xnmos_1p2$$202595372_3v256x8m81_1 pmos_5p04310591302041_3v256x8m81_1/D nmos_5p0431059130208_3v256x8m81_4/D
+ pmos_5p04310591302041_3v256x8m81_1/S vss nmos_1p2$$202595372_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_0 vdd pmos_5p04310591302079_3v256x8m81_0/D vdd nmos_5p0431059130208_3v256x8m81_1/D
+ pmos_5p04310591302014_3v256x8m81
Xpmos_5p04310591302082_3v256x8m81_0 wen pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D
+ pmos_5p04310591302082_3v256x8m81_0/D wen wen vdd wen vdd wen vdd vdd wen vdd pmos_5p04310591302082_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_1 nmos_5p0431059130208_3v256x8m81_3/D clk vdd vdd
+ pmos_5p04310591302014_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_2 vdd pmos_5p04310591302041_3v256x8m81_1/S vdd pmos_5p04310591302014_3v256x8m81_2/S
+ pmos_5p04310591302014_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_3 vdd wen vdd nmos_5p0431059130208_3v256x8m81_2/S
+ pmos_5p04310591302014_3v256x8m81
Xpmos_5p04310591302014_3v256x8m81_4 nmos_5p0431059130208_3v256x8m81_4/D nmos_5p0431059130208_3v256x8m81_3/D
+ vdd vdd pmos_5p04310591302014_3v256x8m81
Xnmos_5p04310591302078_3v256x8m81_0 pmos_5p04310591302082_3v256x8m81_0/D pmos_5p04310591302082_3v256x8m81_0/D
+ vss vss wen wen wen vss nmos_5p04310591302078_3v256x8m81
.ends

.subckt nmos_1p2$$48629804_3v256x8m81 nmos_5p04310591302039_3v256x8m81_0/D nmos_5p04310591302039_3v256x8m81_0/S_uq0
+ a_118_n34# a_n41_n34# nmos_5p04310591302039_3v256x8m81_0/S VSUBS
Xnmos_5p04310591302039_3v256x8m81_0 nmos_5p04310591302039_3v256x8m81_0/D a_n41_n34#
+ a_118_n34# nmos_5p04310591302039_3v256x8m81_0/S_uq0 nmos_5p04310591302039_3v256x8m81_0/S
+ VSUBS nmos_5p04310591302039_3v256x8m81
.ends

.subckt pmos_5p04310591302087_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=4.6552p pd=22.04u as=4.6552p ps=22.04u w=10.58u l=0.28u
.ends

.subckt pmos_1p2$$47815724_3v256x8m81 pmos_5p04310591302087_3v256x8m81_0/D a_n14_n34#
+ pmos_5p04310591302087_3v256x8m81_0/S w_n133_n65#
Xpmos_5p04310591302087_3v256x8m81_0 pmos_5p04310591302087_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302087_3v256x8m81_0/S pmos_5p04310591302087_3v256x8m81
.ends

.subckt nmos_5p04310591302084_3v256x8m81 D_uq2 D_uq1 D_uq0 a_1394_n44# D a_2357_n44#
+ a_1073_n44# a_2036_n44# a_n51_n44# a_1715_n44# a_752_n44# S_uq9 S_uq8 S_uq7 a_n532_n44#
+ S_uq6 S_uq5 a_431_n44# S_uq4 a_1554_n44# a_591_n44# S_uq2 S_uq3 a_2197_n44# S_uq1
+ a_n211_n44# S_uq0 S a_110_n44# a_1876_n44# a_1233_n44# a_270_n44# D_uq8 D_uq7 a_912_n44#
+ D_uq6 a_2518_n44# D_uq4 D_uq5 D_uq3 a_n372_n44# VSUBS
X0 S_uq6 a_270_n44# D_uq6 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X1 D_uq1 a_1715_n44# S_uq2 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.90167p ps=3.96u w=3.435u l=0.28u
X2 D_uq6 a_110_n44# S_uq7 VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X3 D a_2036_n44# S_uq1 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X4 S_uq7 a_n51_n44# D_uq7 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X5 S_uq5 a_591_n44# D_uq5 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X6 D_uq3 a_1073_n44# S_uq4 VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X7 D_uq5 a_431_n44# S_uq6 VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X8 D_uq0 a_2357_n44# S VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X9 D_uq2 a_1394_n44# S_uq3 VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X10 S_uq8 a_n372_n44# D_uq8 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X11 D_uq4 a_752_n44# S_uq5 VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X12 S_uq0 a_2518_n44# D_uq0 VSUBS nfet_03v3 ad=1.5114p pd=7.75u as=0.90167p ps=3.96u w=3.435u l=0.28u
X13 S_uq3 a_1233_n44# D_uq3 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X14 S_uq1 a_1876_n44# D_uq1 VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X15 D_uq7 a_n211_n44# S_uq8 VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X16 S a_2197_n44# D VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=0.90167p ps=3.96u w=3.435u l=0.28u
X17 S_uq2 a_1554_n44# D_uq2 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
X18 D_uq8 a_n532_n44# S_uq9 VSUBS nfet_03v3 ad=0.8931p pd=3.955u as=1.5114p ps=7.75u w=3.435u l=0.28u
X19 S_uq4 a_912_n44# D_uq4 VSUBS nfet_03v3 ad=0.90167p pd=3.96u as=0.8931p ps=3.955u w=3.435u l=0.28u
.ends

.subckt nmos_1p2$$48308268_3v256x8m81 nmos_5p04310591302084_3v256x8m81_0/S_uq5 nmos_5p04310591302084_3v256x8m81_0/a_752_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_1073_n44# nmos_5p04310591302084_3v256x8m81_0/S_uq4
+ nmos_5p04310591302084_3v256x8m81_0/D nmos_5p04310591302084_3v256x8m81_0/a_2036_n44#
+ nmos_5p04310591302084_3v256x8m81_0/S_uq3 nmos_5p04310591302084_3v256x8m81_0/S_uq2
+ nmos_5p04310591302084_3v256x8m81_0/S_uq1 nmos_5p04310591302084_3v256x8m81_0/S_uq0
+ nmos_5p04310591302084_3v256x8m81_0/a_431_n44# nmos_5p04310591302084_3v256x8m81_0/a_1715_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_591_n44# nmos_5p04310591302084_3v256x8m81_0/a_n532_n44#
+ nmos_5p04310591302084_3v256x8m81_0/D_uq8 nmos_5p04310591302084_3v256x8m81_0/D_uq7
+ nmos_5p04310591302084_3v256x8m81_0/a_110_n44# nmos_5p04310591302084_3v256x8m81_0/D_uq6
+ nmos_5p04310591302084_3v256x8m81_0/a_270_n44# nmos_5p04310591302084_3v256x8m81_0/a_1554_n44#
+ nmos_5p04310591302084_3v256x8m81_0/D_uq5 nmos_5p04310591302084_3v256x8m81_0/a_2197_n44#
+ nmos_5p04310591302084_3v256x8m81_0/D_uq4 nmos_5p04310591302084_3v256x8m81_0/a_n211_n44#
+ nmos_5p04310591302084_3v256x8m81_0/D_uq3 nmos_5p04310591302084_3v256x8m81_0/D_uq2
+ nmos_5p04310591302084_3v256x8m81_0/D_uq1 nmos_5p04310591302084_3v256x8m81_0/D_uq0
+ nmos_5p04310591302084_3v256x8m81_0/a_912_n44# nmos_5p04310591302084_3v256x8m81_0/a_1233_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_1876_n44# nmos_5p04310591302084_3v256x8m81_0/S
+ nmos_5p04310591302084_3v256x8m81_0/a_2518_n44# nmos_5p04310591302084_3v256x8m81_0/a_n372_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_1394_n44# nmos_5p04310591302084_3v256x8m81_0/a_2357_n44#
+ nmos_5p04310591302084_3v256x8m81_0/S_uq9 nmos_5p04310591302084_3v256x8m81_0/S_uq8
+ nmos_5p04310591302084_3v256x8m81_0/a_n51_n44# nmos_5p04310591302084_3v256x8m81_0/S_uq7
+ VSUBS nmos_5p04310591302084_3v256x8m81_0/S_uq6
Xnmos_5p04310591302084_3v256x8m81_0 nmos_5p04310591302084_3v256x8m81_0/D_uq2 nmos_5p04310591302084_3v256x8m81_0/D_uq1
+ nmos_5p04310591302084_3v256x8m81_0/D_uq0 nmos_5p04310591302084_3v256x8m81_0/a_1394_n44#
+ nmos_5p04310591302084_3v256x8m81_0/D nmos_5p04310591302084_3v256x8m81_0/a_2357_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_1073_n44# nmos_5p04310591302084_3v256x8m81_0/a_2036_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_n51_n44# nmos_5p04310591302084_3v256x8m81_0/a_1715_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_752_n44# nmos_5p04310591302084_3v256x8m81_0/S_uq9
+ nmos_5p04310591302084_3v256x8m81_0/S_uq8 nmos_5p04310591302084_3v256x8m81_0/S_uq7
+ nmos_5p04310591302084_3v256x8m81_0/a_n532_n44# nmos_5p04310591302084_3v256x8m81_0/S_uq6
+ nmos_5p04310591302084_3v256x8m81_0/S_uq5 nmos_5p04310591302084_3v256x8m81_0/a_431_n44#
+ nmos_5p04310591302084_3v256x8m81_0/S_uq4 nmos_5p04310591302084_3v256x8m81_0/a_1554_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_591_n44# nmos_5p04310591302084_3v256x8m81_0/S_uq2
+ nmos_5p04310591302084_3v256x8m81_0/S_uq3 nmos_5p04310591302084_3v256x8m81_0/a_2197_n44#
+ nmos_5p04310591302084_3v256x8m81_0/S_uq1 nmos_5p04310591302084_3v256x8m81_0/a_n211_n44#
+ nmos_5p04310591302084_3v256x8m81_0/S_uq0 nmos_5p04310591302084_3v256x8m81_0/S nmos_5p04310591302084_3v256x8m81_0/a_110_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_1876_n44# nmos_5p04310591302084_3v256x8m81_0/a_1233_n44#
+ nmos_5p04310591302084_3v256x8m81_0/a_270_n44# nmos_5p04310591302084_3v256x8m81_0/D_uq8
+ nmos_5p04310591302084_3v256x8m81_0/D_uq7 nmos_5p04310591302084_3v256x8m81_0/a_912_n44#
+ nmos_5p04310591302084_3v256x8m81_0/D_uq6 nmos_5p04310591302084_3v256x8m81_0/a_2518_n44#
+ nmos_5p04310591302084_3v256x8m81_0/D_uq4 nmos_5p04310591302084_3v256x8m81_0/D_uq5
+ nmos_5p04310591302084_3v256x8m81_0/D_uq3 nmos_5p04310591302084_3v256x8m81_0/a_n372_n44#
+ VSUBS nmos_5p04310591302084_3v256x8m81
.ends

.subckt nmos_5p04310591302093_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1576p pd=1.64u as=0.1576p ps=1.64u w=0.28u l=0.56u
.ends

.subckt pmos_1p2$$47330348_3v256x8m81 pmos_5p04310591302041_3v256x8m81_0/D a_n14_89#
+ pmos_5p04310591302041_3v256x8m81_0/S w_n133_n65#
Xpmos_5p04310591302041_3v256x8m81_0 pmos_5p04310591302041_3v256x8m81_0/D a_n14_89#
+ w_n133_n65# pmos_5p04310591302041_3v256x8m81_0/S pmos_5p04310591302041_3v256x8m81
.ends

.subckt pmos_5p04310591302089_3v256x8m81 D_uq2 D_uq1 a_2502_n44# D_uq0 a_1699_n44#
+ D a_n67_n44# a_2341_n44# a_1378_n44# a_2020_n44# a_1057_n44# a_n548_n44# S_uq9 S_uq8
+ S_uq7 S_uq6 a_94_n44# S_uq5 a_736_n44# a_n227_n44# S_uq4 S_uq2 S_uq3 a_896_n44#
+ S_uq1 S_uq0 w_n722_n86# S a_415_n44# a_2181_n44# a_1538_n44# a_575_n44# a_1860_n44#
+ D_uq8 D_uq7 a_1217_n44# a_n388_n44# D_uq6 a_254_n44# D_uq4 D_uq5 D_uq3
X0 D_uq8 a_n548_n44# S_uq9 w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=3.7708p ps=18.02u w=8.57u l=0.28u
X1 S_uq5 a_575_n44# D_uq5 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X2 D_uq5 a_415_n44# S_uq6 w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X3 D_uq3 a_1057_n44# S_uq4 w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X4 D a_2020_n44# S_uq1 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X5 S_uq4 a_896_n44# D_uq4 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X6 D_uq4 a_736_n44# S_uq5 w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X7 D_uq2 a_1378_n44# S_uq3 w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X8 D_uq0 a_2341_n44# S w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X9 S_uq7 a_n67_n44# D_uq7 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X10 D_uq1 a_1699_n44# S_uq2 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.24962p ps=9.095u w=8.57u l=0.28u
X11 S_uq0 a_2502_n44# D_uq0 w_n722_n86# pfet_03v3 ad=3.7708p pd=18.02u as=2.24962p ps=9.095u w=8.57u l=0.28u
X12 S_uq8 a_n388_n44# D_uq8 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X13 S_uq3 a_1217_n44# D_uq3 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X14 S_uq1 a_1860_n44# D_uq1 w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X15 S_uq2 a_1538_n44# D_uq2 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
X16 S a_2181_n44# D w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X17 D_uq6 a_94_n44# S_uq7 w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X18 D_uq7 a_n227_n44# S_uq8 w_n722_n86# pfet_03v3 ad=2.2282p pd=9.09u as=2.24962p ps=9.095u w=8.57u l=0.28u
X19 S_uq6 a_254_n44# D_uq6 w_n722_n86# pfet_03v3 ad=2.24962p pd=9.095u as=2.2282p ps=9.09u w=8.57u l=0.28u
.ends

.subckt pmos_5p04310591302073_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.4563p pd=2.275u as=0.7722p ps=4.39u w=1.755u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.7722p pd=4.39u as=0.4563p ps=2.275u w=1.755u l=0.28u
.ends

.subckt pmos_1p2$$48623660_3v256x8m81 a_n42_n34# w_n133_n66# pmos_5p04310591302073_3v256x8m81_0/S_uq0
+ pmos_5p04310591302073_3v256x8m81_0/D a_118_n34# pmos_5p04310591302073_3v256x8m81_0/S
Xpmos_5p04310591302073_3v256x8m81_0 pmos_5p04310591302073_3v256x8m81_0/D a_n42_n34#
+ a_118_n34# w_n133_n66# pmos_5p04310591302073_3v256x8m81_0/S_uq0 pmos_5p04310591302073_3v256x8m81_0/S
+ pmos_5p04310591302073_3v256x8m81
.ends

.subckt pmos_5p04310591302092_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.1848p pd=1.72u as=0.1848p ps=1.72u w=0.42u l=0.465u
.ends

.subckt pmos_5p04310591302091_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=4.004p pd=19.08u as=4.004p ps=19.08u w=9.1u l=0.28u
.ends

.subckt pmos_1p2$$48624684_3v256x8m81 pmos_5p04310591302091_3v256x8m81_0/D a_n14_n34#
+ pmos_5p04310591302091_3v256x8m81_0/S w_n133_n65#
Xpmos_5p04310591302091_3v256x8m81_0 pmos_5p04310591302091_3v256x8m81_0/D a_n14_n34#
+ w_n133_n65# pmos_5p04310591302091_3v256x8m81_0/S pmos_5p04310591302091_3v256x8m81
.ends

.subckt nmos_5p04310591302083_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1646p pd=1.64u as=0.1646p ps=1.64u w=0.35u l=0.28u
.ends

.subckt nmos_5p04310591302090_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1576p pd=1.64u as=0.1576p ps=1.64u w=0.28u l=0.465u
.ends

.subckt pmos_5p04310591302074_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.1848p pd=1.72u as=0.1848p ps=1.72u w=0.42u l=0.56u
.ends

.subckt nmos_5p04310591302085_3v256x8m81 D_uq1 D_uq0 a_530_n44# D a_n112_n44# a_209_n44#
+ a_369_n44# a_48_n44# S_uq1 S_uq0 S VSUBS
X0 D_uq1 a_n112_n44# S_uq1 VSUBS nfet_03v3 ad=1.2103p pd=5.175u as=2.0482p ps=10.19u w=4.655u l=0.28u
X1 S_uq0 a_369_n44# D VSUBS nfet_03v3 ad=1.22192p pd=5.18u as=1.2103p ps=5.175u w=4.655u l=0.28u
X2 D a_209_n44# S VSUBS nfet_03v3 ad=1.2103p pd=5.175u as=1.22192p ps=5.18u w=4.655u l=0.28u
X3 D_uq0 a_530_n44# S_uq0 VSUBS nfet_03v3 ad=2.0482p pd=10.19u as=1.22192p ps=5.18u w=4.655u l=0.28u
X4 S a_48_n44# D_uq1 VSUBS nfet_03v3 ad=1.22192p pd=5.18u as=1.2103p ps=5.175u w=4.655u l=0.28u
.ends

.subckt nmos_1p2$$48306220_3v256x8m81 a_195_n34# a_n125_n34# a_355_n34# nmos_5p04310591302085_3v256x8m81_0/S_uq1
+ nmos_5p04310591302085_3v256x8m81_0/S_uq0 a_34_n34# nmos_5p04310591302085_3v256x8m81_0/D
+ nmos_5p04310591302085_3v256x8m81_0/D_uq1 nmos_5p04310591302085_3v256x8m81_0/D_uq0
+ nmos_5p04310591302085_3v256x8m81_0/S VSUBS a_516_n34#
Xnmos_5p04310591302085_3v256x8m81_0 nmos_5p04310591302085_3v256x8m81_0/D_uq1 nmos_5p04310591302085_3v256x8m81_0/D_uq0
+ a_516_n34# nmos_5p04310591302085_3v256x8m81_0/D a_n125_n34# a_195_n34# a_355_n34#
+ a_34_n34# nmos_5p04310591302085_3v256x8m81_0/S_uq1 nmos_5p04310591302085_3v256x8m81_0/S_uq0
+ nmos_5p04310591302085_3v256x8m81_0/S VSUBS nmos_5p04310591302085_3v256x8m81
.ends

.subckt pmos_5p04310591302094_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.3872p pd=2.64u as=0.3872p ps=2.64u w=0.88u l=0.28u
.ends

.subckt nmos_5p04310591302086_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.6182p pd=3.69u as=0.6182p ps=3.69u w=1.405u l=0.28u
.ends

.subckt nmos_1p2$$48302124_3v256x8m81 nmos_5p04310591302086_3v256x8m81_0/S a_n14_n34#
+ nmos_5p04310591302086_3v256x8m81_0/D VSUBS
Xnmos_5p04310591302086_3v256x8m81_0 nmos_5p04310591302086_3v256x8m81_0/D a_n14_n34#
+ nmos_5p04310591302086_3v256x8m81_0/S VSUBS nmos_5p04310591302086_3v256x8m81
.ends

.subckt gen_3v256x8_3v256x8m81 tblhl IGWEN cen clk WEN GWE VDD_uq3 pmos_5p04310591302088_3v256x8m81_0/D
+ men VSS wen_v2_3v256x8m81_0/wen VDD_uq2 VDD
Xpmos_5p04310591302088_3v256x8m81_0 pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ VDD_uq3 VDD_uq3 VDD_uq3 VDD_uq3 VDD_uq3 pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ VDD_uq3 VDD_uq3 pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_5p04310591302088_3v256x8m81
Xwen_v2_3v256x8m81_0 clk wen_v2_3v256x8m81_0/wen GWE VDD IGWEN VSS wen_v2_3v256x8m81
Xnmos_1p2$$48629804_3v256x8m81_0 pmos_5p04310591302051_3v256x8m81_0/D VSS nmos_1p2$$46563372_3v256x8m81_2/nmos_5p0431059130208_3v256x8m81_0/S
+ nmos_1p2$$46563372_3v256x8m81_2/nmos_5p0431059130208_3v256x8m81_0/S VSS VSS nmos_1p2$$48629804_3v256x8m81
Xpmos_1p2$$47815724_3v256x8m81_0 VDD_uq2 tblhl pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S
+ VDD_uq2 pmos_1p2$$47815724_3v256x8m81
Xpmos_1p2$$47815724_3v256x8m81_1 pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S VDD_uq2 VDD_uq2
+ pmos_1p2$$47815724_3v256x8m81
Xnmos_1p2$$48308268_3v256x8m81_0 VSS pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ VSS men pmos_5p04310591302088_3v256x8m81_0/D VSS VSS VSS VSS pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ men men pmos_5p04310591302088_3v256x8m81_0/D men pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D men pmos_5p04310591302088_3v256x8m81_0/D men
+ pmos_5p04310591302088_3v256x8m81_0/D men men men men pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D VSS pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ VSS VSS pmos_5p04310591302088_3v256x8m81_0/D VSS VSS VSS nmos_1p2$$48308268_3v256x8m81
Xpmos_1p2$$47815724_3v256x8m81_2 pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S
+ tblhl VDD_uq2 VDD_uq2 pmos_1p2$$47815724_3v256x8m81
Xnmos_5p04310591302093_3v256x8m81_0 pmos_5p04310591302074_3v256x8m81_0/D clk VSS VSS
+ nmos_5p04310591302093_3v256x8m81
Xnmos_5p04310591302093_3v256x8m81_1 pmos_5p04310591302074_3v256x8m81_1/D pmos_5p04310591302074_3v256x8m81_0/D
+ VSS VSS nmos_5p04310591302093_3v256x8m81
Xpmos_1p2$$47815724_3v256x8m81_3 VDD_uq2 pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S VDD_uq2 pmos_1p2$$47815724_3v256x8m81
Xpmos_1p2$$47330348_3v256x8m81_0 pmos_1p2$$46273580_3v256x8m81_0/pmos_5p0431059130203_3v256x8m81_0/D
+ nmos_1p2$$47342636_3v256x8m81_1/nmos_5p04310591302053_3v256x8m81_0/S nmos_1p2$$46563372_3v256x8m81_2/nmos_5p0431059130208_3v256x8m81_0/S
+ VDD_uq2 pmos_1p2$$47330348_3v256x8m81
Xpmos_5p04310591302089_3v256x8m81_0 men men pmos_5p04310591302088_3v256x8m81_0/D men
+ pmos_5p04310591302088_3v256x8m81_0/D men pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D VDD_uq3 VDD_uq3 VDD_uq3 VDD_uq3 pmos_5p04310591302088_3v256x8m81_0/D
+ VDD_uq3 pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ VDD_uq3 VDD_uq3 VDD_uq3 pmos_5p04310591302088_3v256x8m81_0/D VDD_uq3 VDD_uq3 VDD_uq3
+ VDD_uq3 pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ men men pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D
+ men pmos_5p04310591302088_3v256x8m81_0/D men men men pmos_5p04310591302089_3v256x8m81
Xpmos_1p2$$48623660_3v256x8m81_0 pmos_5p04310591302094_3v256x8m81_0/D VDD VDD pmos_1p2$$48623660_3v256x8m81_0/pmos_5p04310591302073_3v256x8m81_0/D
+ pmos_5p04310591302094_3v256x8m81_0/D VDD pmos_1p2$$48623660_3v256x8m81
Xpmos_1p2$$47815724_3v256x8m81_4 pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S VDD_uq2 VDD_uq2
+ pmos_1p2$$47815724_3v256x8m81
Xpmos_1p2$$47815724_3v256x8m81_5 pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$48624684_3v256x8m81_2/pmos_5p04310591302091_3v256x8m81_0/S VDD_uq2 VDD_uq2
+ pmos_1p2$$47815724_3v256x8m81
Xpmos_1p2$$47815724_3v256x8m81_6 VDD_uq2 pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S VDD_uq2 pmos_1p2$$47815724_3v256x8m81
Xpmos_1p2$$47815724_3v256x8m81_7 VDD_uq2 pmos_1p2$$48624684_3v256x8m81_2/pmos_5p04310591302091_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S VDD_uq2 pmos_1p2$$47815724_3v256x8m81
Xnmos_1p2$$47342636_3v256x8m81_0 nmos_1p2$$47342636_3v256x8m81_1/nmos_5p04310591302053_3v256x8m81_0/S
+ clk VSS VSS nmos_1p2$$47342636_3v256x8m81
Xpmos_5p04310591302092_3v256x8m81_0 pmos_5p04310591302092_3v256x8m81_0/D pmos_5p04310591302074_3v256x8m81_1/D
+ VDD VDD pmos_5p04310591302092_3v256x8m81
Xnmos_1p2$$47342636_3v256x8m81_1 VSS men VSS nmos_1p2$$47342636_3v256x8m81_1/nmos_5p04310591302053_3v256x8m81_0/S
+ nmos_1p2$$47342636_3v256x8m81
Xpmos_1p2$$48624684_3v256x8m81_0 pmos_1p2$$48624684_3v256x8m81_2/pmos_5p04310591302091_3v256x8m81_0/S
+ pmos_5p04310591302051_3v256x8m81_0/D VDD_uq2 VDD_uq2 pmos_1p2$$48624684_3v256x8m81
Xpmos_1p2$$48624684_3v256x8m81_1 pmos_1p2$$48624684_3v256x8m81_2/pmos_5p04310591302091_3v256x8m81_0/S
+ pmos_1p2$$48623660_3v256x8m81_0/pmos_5p04310591302073_3v256x8m81_0/D VDD_uq2 VDD_uq2
+ pmos_1p2$$48624684_3v256x8m81
Xpmos_1p2$$46273580_3v256x8m81_0 VDD_uq2 pmos_5p04310591302051_3v256x8m81_0/D VDD_uq2
+ VDD_uq2 pmos_5p04310591302051_3v256x8m81_0/D pmos_1p2$$46273580_3v256x8m81_0/pmos_5p0431059130203_3v256x8m81_0/D
+ pmos_1p2$$46273580_3v256x8m81
Xpmos_1p2$$48624684_3v256x8m81_2 VDD_uq2 clk pmos_1p2$$48624684_3v256x8m81_2/pmos_5p04310591302091_3v256x8m81_0/S
+ VDD_uq2 pmos_1p2$$48624684_3v256x8m81
Xnmos_5p04310591302083_3v256x8m81_0 pmos_5p04310591302094_3v256x8m81_0/D pmos_5p04310591302092_3v256x8m81_0/D
+ VSS VSS nmos_5p04310591302083_3v256x8m81
Xnmos_5p04310591302090_3v256x8m81_0 pmos_5p04310591302092_3v256x8m81_0/D pmos_5p04310591302074_3v256x8m81_1/D
+ VSS VSS nmos_5p04310591302090_3v256x8m81
Xpmos_5p04310591302074_3v256x8m81_0 pmos_5p04310591302074_3v256x8m81_0/D clk VDD VDD
+ pmos_5p04310591302074_3v256x8m81
Xpmos_5p04310591302074_3v256x8m81_1 pmos_5p04310591302074_3v256x8m81_1/D pmos_5p04310591302074_3v256x8m81_0/D
+ VDD VDD pmos_5p04310591302074_3v256x8m81
Xnmos_1p2$$48306220_3v256x8m81_0 pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S
+ VSS VSS pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S pmos_5p04310591302088_3v256x8m81_0/D
+ pmos_5p04310591302088_3v256x8m81_0/D pmos_5p04310591302088_3v256x8m81_0/D VSS VSS
+ pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S nmos_1p2$$48306220_3v256x8m81
Xpmos_5p04310591302051_3v256x8m81_0 pmos_5p04310591302051_3v256x8m81_0/D nmos_1p2$$46563372_3v256x8m81_2/nmos_5p0431059130208_3v256x8m81_0/S
+ nmos_1p2$$46563372_3v256x8m81_2/nmos_5p0431059130208_3v256x8m81_0/S VDD_uq2 VDD_uq2
+ VDD_uq2 pmos_5p04310591302051_3v256x8m81
Xnmos_1p2$$46563372_3v256x8m81_0 nmos_1p2$$46563372_3v256x8m81_0/nmos_5p0431059130208_3v256x8m81_0/D
+ nmos_1p2$$47342636_3v256x8m81_1/nmos_5p04310591302053_3v256x8m81_0/S VSS VSS nmos_1p2$$46563372_3v256x8m81
Xpmos_5p04310591302094_3v256x8m81_0 pmos_5p04310591302094_3v256x8m81_0/D pmos_5p04310591302092_3v256x8m81_0/D
+ VDD VDD pmos_5p04310591302094_3v256x8m81
Xnmos_1p2$$46563372_3v256x8m81_1 VSS pmos_5p04310591302051_3v256x8m81_0/D pmos_1p2$$46273580_3v256x8m81_0/pmos_5p0431059130203_3v256x8m81_0/D
+ VSS nmos_1p2$$46563372_3v256x8m81
Xpmos_1p2$$46285868_3v256x8m81_0 VDD_uq2 VDD_uq2 nmos_1p2$$46563372_3v256x8m81_0/nmos_5p0431059130208_3v256x8m81_0/D
+ nmos_1p2$$47342636_3v256x8m81_1/nmos_5p04310591302053_3v256x8m81_0/S pmos_1p2$$46285868_3v256x8m81
Xnmos_1p2$$46551084_3v256x8m81_0 cen nmos_1p2$$47342636_3v256x8m81_1/nmos_5p04310591302053_3v256x8m81_0/S
+ nmos_1p2$$46563372_3v256x8m81_2/nmos_5p0431059130208_3v256x8m81_0/S VSS nmos_1p2$$46551084_3v256x8m81
Xnmos_1p2$$46563372_3v256x8m81_2 pmos_1p2$$46273580_3v256x8m81_0/pmos_5p0431059130203_3v256x8m81_0/D
+ nmos_1p2$$46563372_3v256x8m81_0/nmos_5p0431059130208_3v256x8m81_0/D nmos_1p2$$46563372_3v256x8m81_2/nmos_5p0431059130208_3v256x8m81_0/S
+ VSS nmos_1p2$$46563372_3v256x8m81
Xpmos_1p2$$46285868_3v256x8m81_1 VDD_uq2 nmos_1p2$$46563372_3v256x8m81_2/nmos_5p0431059130208_3v256x8m81_0/S
+ cen nmos_1p2$$46563372_3v256x8m81_0/nmos_5p0431059130208_3v256x8m81_0/D pmos_1p2$$46285868_3v256x8m81
Xnmos_1p2$$48302124_3v256x8m81_0 VSS pmos_5p04310591302094_3v256x8m81_0/D pmos_1p2$$48623660_3v256x8m81_0/pmos_5p04310591302073_3v256x8m81_0/D
+ VSS nmos_1p2$$48302124_3v256x8m81
X0 a_8790_2243# tblhl pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S VSS nfet_03v3 ad=0.5499p pd=2.635u as=0.5499p ps=2.635u w=2.115u l=0.28u
X1 a_3606_4291# men VDD_uq2 VDD_uq2 pfet_03v3 ad=0.2769p pd=1.585u as=0.50587p ps=3.08u w=1.065u l=0.28u
X2 a_7891_338# pmos_1p2$$48624684_3v256x8m81_2/pmos_5p04310591302091_3v256x8m81_0/S pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S VSS nfet_03v3 ad=2.2009p pd=8.985u as=2.2009p ps=8.985u w=8.465u l=0.28u
X3 a_6888_183# clk a_6728_183# VSS nfet_03v3 ad=2.7521p pd=11.105u as=2.7521p ps=11.105u w=10.585u l=0.28u
X4 VSS pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S a_7891_338# VSS nfet_03v3 ad=3.93622p pd=17.86u as=2.2009p ps=8.985u w=8.465u l=0.28u
X5 pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S tblhl a_8470_2243# VSS nfet_03v3 ad=0.5499p pd=2.635u as=0.5499p ps=2.635u w=2.115u l=0.28u
X6 a_8470_2243# pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S VSS VSS nfet_03v3 ad=0.5499p pd=2.635u as=0.96232p ps=5.14u w=2.115u l=0.28u
X7 pmos_1p2$$48624684_3v256x8m81_2/pmos_5p04310591302091_3v256x8m81_0/S pmos_5p04310591302051_3v256x8m81_0/D a_6888_183# VSS nfet_03v3 ad=5.2925p pd=22.17u as=2.7521p ps=11.105u w=10.585u l=0.28u
X8 a_7571_338# pmos_1p2$$47815724_3v256x8m81_3/pmos_5p04310591302087_3v256x8m81_0/S VSS VSS nfet_03v3 ad=2.2009p pd=8.985u as=3.85157p ps=17.84u w=8.465u l=0.28u
X9 pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S pmos_1p2$$48624684_3v256x8m81_2/pmos_5p04310591302091_3v256x8m81_0/S a_7571_338# VSS nfet_03v3 ad=2.2009p pd=8.985u as=2.2009p ps=8.985u w=8.465u l=0.28u
X10 a_6728_183# pmos_1p2$$48623660_3v256x8m81_0/pmos_5p04310591302073_3v256x8m81_0/D VSS VSS nfet_03v3 ad=2.7521p pd=11.105u as=4.6574p ps=22.05u w=10.585u l=0.28u
X11 nmos_1p2$$47342636_3v256x8m81_1/nmos_5p04310591302053_3v256x8m81_0/S clk a_3606_4291# VDD_uq2 pfet_03v3 ad=0.50587p pd=3.08u as=0.2769p ps=1.585u w=1.065u l=0.28u
X12 VSS pmos_1p2$$47815724_3v256x8m81_7/pmos_5p04310591302087_3v256x8m81_0/S a_8790_2243# VSS nfet_03v3 ad=0.99405p pd=5.17u as=0.5499p ps=2.635u w=2.115u l=0.28u
.ends

.subckt control_3v256x8_3v256x8m81 VDD RYS[7] RYS[6] RYS[5] RYS[4] RYS[3] RYS[2] RYS[1]
+ RYS[0] LYS[0] LYS[1] LYS[2] LYS[3] LYS[6] LYS[5] LYS[4] LYS[7] tblhl IGWEN xb[3]
+ xb[2] xb[0] xa[7] xa[6] xa[5] xa[4] xa[2] A[0] xb[1] xc[3] xc[1] xc[2] xa[1] A[9]
+ A[7] CLK A[2] A[1] A[6] A[3] A[4] A[5] A[8] GWE GWEN VSS_uq2 VSS_uq5 VDD_uq0 VDD_uq5
+ ypredec1_3v256x8m81_0/ly[1] ypredec1_3v256x8m81_0/ly[2] men VDD_uq4 ypredec1_3v256x8m81_0/ly[4]
+ xa[3] ypredec1_3v256x8m81_0/ly[5] ypredec1_3v256x8m81_0/ly[6] xa[0] ypredec1_3v256x8m81_0/ly[7]
+ CEN prexdec_top_3v256x8m81_0/xpredec0_3v256x8m81_1/vdd VDD_uq1 VDD_uq2 xc[0] prexdec_top_3v256x8m81_0/xpredec1_3v256x8m81_0/xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd
+ VDD_uq6 VSS gen_3v256x8_3v256x8m81_0/VDD_uq2 VDD_uq3
Xypredec1_3v256x8m81_0 ypredec1_3v256x8m81_0/ly[5] ypredec1_3v256x8m81_0/ly[4] ypredec1_3v256x8m81_0/ly[7]
+ ypredec1_3v256x8m81_0/ly[2] ypredec1_3v256x8m81_0/ly[1] LYS[7] RYS[0] RYS[1] RYS[2]
+ RYS[3] RYS[4] RYS[5] RYS[6] RYS[7] ypredec1_3v256x8m81_0/ly[6] men A[0] A[1] A[2]
+ CLK A[1] VDD_uq4 A[0] VDD A[2] VDD VDD_uq6 VSS VDD_uq1 VDD_uq2 ypredec1_3v256x8m81
Xprexdec_top_3v256x8m81_0 A[5] A[9] xb[3] xc[1] xc[2] xc[3] xb[1] xb[2] xb[0] xa[1]
+ xa[2] xa[4] xa[5] xa[6] xa[7] A[3] A[6] A[8] A[4] xa[0] VSS xa[3] CLK VSS VSS VDD_uq3
+ VSS VDD_uq3 A[7] xc[0] men prexdec_top_3v256x8m81_0/xpredec0_3v256x8m81_1/vdd prexdec_top_3v256x8m81_0/xpredec1_3v256x8m81_0/xpredec1_bot_3v256x8m81_2/alatch_3v256x8m81_0/vdd
+ CLK VDD_uq3 VSS prexdec_top_3v256x8m81
Xgen_3v256x8_3v256x8m81_0 tblhl IGWEN CEN CLK gen_3v256x8_3v256x8m81_0/WEN GWE VDD_uq6
+ gen_3v256x8_3v256x8m81_0/pmos_5p04310591302088_3v256x8m81_0/D men VSS GWEN gen_3v256x8_3v256x8m81_0/VDD_uq2
+ VDD gen_3v256x8_3v256x8m81
.ends

.subckt pmos_5p043105913020101_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=1.353p pd=7.03u as=1.353p ps=7.03u w=3.075u l=0.28u
.ends

.subckt nmos_5p043105913020107_3v256x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.6058p pd=2.85u as=1.0252p ps=5.54u w=2.33u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=1.0252p pd=5.54u as=0.6058p ps=2.85u w=2.33u l=0.28u
.ends

.subckt pmos_5p043105913020103_3v256x8m81 D_uq0 D a_265_n44# S_uq0 S a_n56_n44# a_104_n44#
+ w_n230_n86#
X0 D_uq0 a_265_n44# S_uq0 w_n230_n86# pfet_03v3 ad=2.0526p pd=10.21u as=1.22455p ps=5.19u w=4.665u l=0.28u
X1 D a_n56_n44# S w_n230_n86# pfet_03v3 ad=1.2129p pd=5.185u as=2.0526p ps=10.21u w=4.665u l=0.28u
X2 S_uq0 a_104_n44# D w_n230_n86# pfet_03v3 ad=1.22455p pd=5.19u as=1.2129p ps=5.185u w=4.665u l=0.28u
.ends

.subckt pmos_1p2_03_R270_3v256x8m81 a_n69_n138# pmos_5p043105913020103_3v256x8m81_0/S_uq0
+ pmos_5p043105913020103_3v256x8m81_0/S a_90_n138# w_n138_n63# pmos_5p043105913020103_3v256x8m81_0/D_uq0
+ a_251_n138# pmos_5p043105913020103_3v256x8m81_0/D
Xpmos_5p043105913020103_3v256x8m81_0 pmos_5p043105913020103_3v256x8m81_0/D_uq0 pmos_5p043105913020103_3v256x8m81_0/D
+ a_251_n138# pmos_5p043105913020103_3v256x8m81_0/S_uq0 pmos_5p043105913020103_3v256x8m81_0/S
+ a_n69_n138# a_90_n138# w_n138_n63# pmos_5p043105913020103_3v256x8m81
.ends

.subckt pmos_5p043105913020108_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.6669p pd=3.085u as=1.1286p ps=6.01u w=2.565u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=1.1286p pd=6.01u as=0.6669p ps=3.085u w=2.565u l=0.28u
.ends

.subckt pmos_1p2_01_R270_3v256x8m81 pmos_5p043105913020108_3v256x8m81_0/S_uq0 pmos_5p043105913020108_3v256x8m81_0/D
+ w_n246_n93# a_118_n33# pmos_5p043105913020108_3v256x8m81_0/S a_n41_n33#
Xpmos_5p043105913020108_3v256x8m81_0 pmos_5p043105913020108_3v256x8m81_0/D a_n41_n33#
+ a_118_n33# w_n246_n93# pmos_5p043105913020108_3v256x8m81_0/S_uq0 pmos_5p043105913020108_3v256x8m81_0/S
+ pmos_5p043105913020108_3v256x8m81
.ends

.subckt nmos_1p2_02_R270_3v256x8m81 nmos_5p04310591302044_3v256x8m81_0/S a_n14_n33#
+ nmos_5p04310591302044_3v256x8m81_0/D VSUBS
Xnmos_5p04310591302044_3v256x8m81_0 nmos_5p04310591302044_3v256x8m81_0/D a_n14_n33#
+ nmos_5p04310591302044_3v256x8m81_0/S VSUBS nmos_5p04310591302044_3v256x8m81
.ends

.subckt nmos_5p043105913020109_3v256x8m81 D a_n28_n44# a_132_n44# S_uq0 S VSUBS
X0 D a_n28_n44# S VSUBS nfet_03v3 ad=0.4004p pd=2.06u as=0.6776p ps=3.96u w=1.54u l=0.28u
X1 S_uq0 a_132_n44# D VSUBS nfet_03v3 ad=0.6776p pd=3.96u as=0.4004p ps=2.06u w=1.54u l=0.28u
.ends

.subckt pmos_5p043105913020110_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.3256p pd=2.36u as=0.3256p ps=2.36u w=0.74u l=0.28u
.ends

.subckt pmos_5p043105913020104_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=0.4004p pd=2.06u as=0.6776p ps=3.96u w=1.54u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=0.6776p pd=3.96u as=0.4004p ps=2.06u w=1.54u l=0.28u
.ends

.subckt pmos_1p2_02_R270_3v256x8m81 a_118_n33# a_n41_n33# pmos_5p043105913020104_3v256x8m81_0/D
+ w_n138_n63# pmos_5p043105913020104_3v256x8m81_0/S_uq0 pmos_5p043105913020104_3v256x8m81_0/S
Xpmos_5p043105913020104_3v256x8m81_0 pmos_5p043105913020104_3v256x8m81_0/D a_n41_n33#
+ a_118_n33# w_n138_n63# pmos_5p043105913020104_3v256x8m81_0/S_uq0 pmos_5p043105913020104_3v256x8m81_0/S
+ pmos_5p043105913020104_3v256x8m81
.ends

.subckt nmos_5p043105913020106_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.1601p pd=1.64u as=0.1601p ps=1.64u w=0.305u l=0.28u
.ends

.subckt pmos_5p043105913020105_3v256x8m81 D a_0_n44# w_n174_n86# S
X0 D a_0_n44# S w_n174_n86# pfet_03v3 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.28u
.ends

.subckt xdec_3v256x8m81 RWL LWL men xc xb xa m2_11898_n156# m2_9070_n156# m2_7748_n156#
+ m2_8806_n156# m2_10577_n156# m2_10840_n156# m2_7219_n156# m2_7483_n156# m2_11634_n156#
+ m2_8277_n156# m2_12427_n156# m2_8541_n156# m2_11105_n156# m2_11370_n156# m2_8012_n156#
+ m2_12163_n156# vss vdd
Xnmos_5p043105913020107_3v256x8m81_0 LWL pmos_1p2_01_R270_3v256x8m81_1/pmos_5p043105913020108_3v256x8m81_0/D
+ pmos_1p2_01_R270_3v256x8m81_1/pmos_5p043105913020108_3v256x8m81_0/D vss vss vss
+ nmos_5p043105913020107_3v256x8m81
Xpmos_1p2_03_R270_3v256x8m81_0 pmos_1p2_01_R270_3v256x8m81_1/pmos_5p043105913020108_3v256x8m81_0/D
+ LWL LWL pmos_1p2_01_R270_3v256x8m81_1/pmos_5p043105913020108_3v256x8m81_0/D vdd
+ vdd pmos_1p2_01_R270_3v256x8m81_1/pmos_5p043105913020108_3v256x8m81_0/D vdd pmos_1p2_03_R270_3v256x8m81
Xnmos_5p043105913020107_3v256x8m81_1 RWL pmos_1p2_01_R270_3v256x8m81_0/pmos_5p043105913020108_3v256x8m81_0/D
+ pmos_1p2_01_R270_3v256x8m81_0/pmos_5p043105913020108_3v256x8m81_0/D vss vss vss
+ nmos_5p043105913020107_3v256x8m81
Xpmos_1p2_01_R270_3v256x8m81_0 vdd pmos_1p2_01_R270_3v256x8m81_0/pmos_5p043105913020108_3v256x8m81_0/D
+ vdd nmos_5p043105913020109_3v256x8m81_0/S vdd nmos_5p043105913020109_3v256x8m81_0/S
+ pmos_1p2_01_R270_3v256x8m81
Xpmos_1p2_01_R270_3v256x8m81_1 vdd pmos_1p2_01_R270_3v256x8m81_1/pmos_5p043105913020108_3v256x8m81_0/D
+ vdd nmos_5p043105913020109_3v256x8m81_0/S vdd nmos_5p043105913020109_3v256x8m81_0/S
+ pmos_1p2_01_R270_3v256x8m81
Xnmos_1p2_02_R270_3v256x8m81_0 nmos_5p043105913020109_3v256x8m81_0/S pmos_5p043105913020105_3v256x8m81_3/S
+ vss vss nmos_1p2_02_R270_3v256x8m81
Xnmos_5p043105913020109_3v256x8m81_0 men pmos_5p043105913020110_3v256x8m81_0/S pmos_5p043105913020110_3v256x8m81_0/S
+ nmos_5p043105913020109_3v256x8m81_0/S nmos_5p043105913020109_3v256x8m81_0/S vss
+ nmos_5p043105913020109_3v256x8m81
Xpmos_5p043105913020103_3v256x8m81_0 vdd vdd pmos_1p2_01_R270_3v256x8m81_0/pmos_5p043105913020108_3v256x8m81_0/D
+ RWL RWL pmos_1p2_01_R270_3v256x8m81_0/pmos_5p043105913020108_3v256x8m81_0/D pmos_1p2_01_R270_3v256x8m81_0/pmos_5p043105913020108_3v256x8m81_0/D
+ vdd pmos_5p043105913020103_3v256x8m81
Xpmos_5p043105913020110_3v256x8m81_0 vdd pmos_5p043105913020105_3v256x8m81_3/S vdd
+ pmos_5p043105913020110_3v256x8m81_0/S pmos_5p043105913020110_3v256x8m81
Xpmos_1p2_02_R270_3v256x8m81_0 pmos_5p043105913020105_3v256x8m81_3/S pmos_5p043105913020105_3v256x8m81_3/S
+ men vdd nmos_5p043105913020109_3v256x8m81_0/S nmos_5p043105913020109_3v256x8m81_0/S
+ pmos_1p2_02_R270_3v256x8m81
Xnmos_5p043105913020106_3v256x8m81_0 vss pmos_5p043105913020105_3v256x8m81_3/S pmos_5p043105913020110_3v256x8m81_0/S
+ vss nmos_5p043105913020106_3v256x8m81
Xpmos_5p043105913020105_3v256x8m81_1 pmos_5p043105913020105_3v256x8m81_3/S xb vdd
+ vdd pmos_5p043105913020105_3v256x8m81
Xpmos_5p043105913020105_3v256x8m81_2 vdd xa vdd pmos_5p043105913020105_3v256x8m81_3/S
+ pmos_5p043105913020105_3v256x8m81
Xpmos_5p043105913020105_3v256x8m81_3 vdd xc vdd pmos_5p043105913020105_3v256x8m81_3/S
+ pmos_5p043105913020105_3v256x8m81
X0 vss xc a_9450_422# vss nfet_03v3 ad=0.88935p pd=4.15u as=0.29032p ps=1.865u w=1.47u l=0.28u
X1 vss nmos_5p043105913020109_3v256x8m81_0/S pmos_1p2_01_R270_3v256x8m81_1/pmos_5p043105913020108_3v256x8m81_0/D vss nfet_03v3 ad=0.2796p pd=4.9u as=1.0252p ps=5.54u w=2.33u l=0.28u
X2 a_9450_280# xa pmos_5p043105913020105_3v256x8m81_3/S vss nfet_03v3 ad=0.31605p pd=1.9u as=0.74235p ps=3.95u w=1.47u l=0.28u
X3 a_9450_422# xb a_9450_280# vss nfet_03v3 ad=0.29032p pd=1.865u as=0.31605p ps=1.9u w=1.47u l=0.28u
X4 vss nmos_5p043105913020109_3v256x8m81_0/S pmos_1p2_01_R270_3v256x8m81_0/pmos_5p043105913020108_3v256x8m81_0/D vss nfet_03v3 ad=1.15335p pd=5.65u as=1.0718p ps=5.58u w=2.33u l=0.28u
.ends

.subckt xdec8_3v256x8m81 LWL[5] LWL[4] LWL[2] RWL[5] RWL[4] RWL[2] RWL[7] LWL[1] LWL[7]
+ LWL[6] LWL[0] LWL[3] xb xa[4] xa[7] xa[1] xb_uq3 xb_uq6 xc_uq0 xc_uq2 xc_uq3 xc_uq5
+ xb_uq2 xb_uq0 xa[3] xb_uq5 xa[0] xa[6] xdec_3v256x8m81_7/m2_10577_n156# RWL[3] xc_uq4
+ xc_uq1 xb_uq4 xdec_3v256x8m81_7/m2_7219_n156# xb_uq1 xdec_3v256x8m81_7/m2_11634_n156#
+ xa[5] xa[2] RWL[0] xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_12427_n156#
+ RWL[6] xdec_3v256x8m81_7/m2_11898_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_9070_n156#
+ men xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_8541_n156#
+ xdec_3v256x8m81_7/m2_12163_n156# xdec_3v256x8m81_7/m2_8277_n156# RWL[1] xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_8012_n156# xc vdd vss xdec_3v256x8m81_7/m2_11105_n156# xc_uq6
Xxdec_3v256x8m81_6 RWL[3] LWL[3] men xc_uq2 xb_uq2 xa[3] xdec_3v256x8m81_7/m2_11898_n156#
+ xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_10577_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_7219_n156#
+ xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_11634_n156# xdec_3v256x8m81_7/m2_8277_n156#
+ xdec_3v256x8m81_7/m2_12427_n156# xdec_3v256x8m81_7/m2_8541_n156# xdec_3v256x8m81_7/m2_11105_n156#
+ xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_8012_n156# xdec_3v256x8m81_7/m2_12163_n156#
+ vss vdd xdec_3v256x8m81
Xxdec_3v256x8m81_7 RWL[1] LWL[1] men xc xb xa[1] xdec_3v256x8m81_7/m2_11898_n156#
+ xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_10577_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_7219_n156#
+ xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_11634_n156# xdec_3v256x8m81_7/m2_8277_n156#
+ xdec_3v256x8m81_7/m2_12427_n156# xdec_3v256x8m81_7/m2_8541_n156# xdec_3v256x8m81_7/m2_11105_n156#
+ xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_8012_n156# xdec_3v256x8m81_7/m2_12163_n156#
+ vss vdd xdec_3v256x8m81
Xxdec_3v256x8m81_0 RWL[6] LWL[6] men xc_uq5 xb_uq5 xa[6] xdec_3v256x8m81_7/m2_11898_n156#
+ xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_10577_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_7219_n156#
+ xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_11634_n156# xdec_3v256x8m81_7/m2_8277_n156#
+ xdec_3v256x8m81_7/m2_12427_n156# xdec_3v256x8m81_7/m2_8541_n156# xdec_3v256x8m81_7/m2_11105_n156#
+ xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_8012_n156# xdec_3v256x8m81_7/m2_12163_n156#
+ vss vdd xdec_3v256x8m81
Xxdec_3v256x8m81_1 RWL[4] LWL[4] men xc_uq3 xb_uq3 xa[4] xdec_3v256x8m81_7/m2_11898_n156#
+ xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_10577_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_7219_n156#
+ xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_11634_n156# xdec_3v256x8m81_7/m2_8277_n156#
+ xdec_3v256x8m81_7/m2_12427_n156# xdec_3v256x8m81_7/m2_8541_n156# xdec_3v256x8m81_7/m2_11105_n156#
+ xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_8012_n156# xdec_3v256x8m81_7/m2_12163_n156#
+ vss vdd xdec_3v256x8m81
Xxdec_3v256x8m81_2 RWL[2] LWL[2] men xc_uq1 xb_uq1 xa[2] xdec_3v256x8m81_7/m2_11898_n156#
+ xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_10577_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_7219_n156#
+ xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_11634_n156# xdec_3v256x8m81_7/m2_8277_n156#
+ xdec_3v256x8m81_7/m2_12427_n156# xdec_3v256x8m81_7/m2_8541_n156# xdec_3v256x8m81_7/m2_11105_n156#
+ xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_8012_n156# xdec_3v256x8m81_7/m2_12163_n156#
+ vss vdd xdec_3v256x8m81
Xxdec_3v256x8m81_3 RWL[0] LWL[0] men xc_uq0 xb_uq0 xa[0] xdec_3v256x8m81_7/m2_11898_n156#
+ xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_10577_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_7219_n156#
+ xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_11634_n156# xdec_3v256x8m81_7/m2_8277_n156#
+ xdec_3v256x8m81_7/m2_12427_n156# xdec_3v256x8m81_7/m2_8541_n156# xdec_3v256x8m81_7/m2_11105_n156#
+ xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_8012_n156# xdec_3v256x8m81_7/m2_12163_n156#
+ vss vdd xdec_3v256x8m81
Xxdec_3v256x8m81_4 RWL[7] LWL[7] men xc_uq6 xb_uq6 xa[7] xdec_3v256x8m81_7/m2_11898_n156#
+ xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_10577_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_7219_n156#
+ xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_11634_n156# xdec_3v256x8m81_7/m2_8277_n156#
+ xdec_3v256x8m81_7/m2_12427_n156# xdec_3v256x8m81_7/m2_8541_n156# xdec_3v256x8m81_7/m2_11105_n156#
+ xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_8012_n156# xdec_3v256x8m81_7/m2_12163_n156#
+ vss vdd xdec_3v256x8m81
Xxdec_3v256x8m81_5 RWL[5] LWL[5] men xc_uq4 xb_uq4 xa[5] xdec_3v256x8m81_7/m2_11898_n156#
+ xdec_3v256x8m81_7/m2_9070_n156# xdec_3v256x8m81_7/m2_7748_n156# xdec_3v256x8m81_7/m2_8806_n156#
+ xdec_3v256x8m81_7/m2_10577_n156# xdec_3v256x8m81_7/m2_10840_n156# xdec_3v256x8m81_7/m2_7219_n156#
+ xdec_3v256x8m81_7/m2_7483_n156# xdec_3v256x8m81_7/m2_11634_n156# xdec_3v256x8m81_7/m2_8277_n156#
+ xdec_3v256x8m81_7/m2_12427_n156# xdec_3v256x8m81_7/m2_8541_n156# xdec_3v256x8m81_7/m2_11105_n156#
+ xdec_3v256x8m81_7/m2_11370_n156# xdec_3v256x8m81_7/m2_8012_n156# xdec_3v256x8m81_7/m2_12163_n156#
+ vss vdd xdec_3v256x8m81
.ends

.subckt xdec32_3v256x8m81 LWL[6] LWL[7] RWL[18] RWL[17] RWL[14] RWL[13] LWL[9] LWL[8]
+ LWL[0] LWL[1] LWL[2] LWL[3] LWL[4] LWL[5] RWL[11] RWL[10] RWL[8] RWL[5] RWL[3] RWL[0]
+ RWL[2] LWL[18] LWL[17] LWL[16] LWL[15] LWL[14] LWL[13] LWL[12] LWL[11] LWL[10] RWL[6]
+ LWL[28] LWL[27] LWL[26] LWL[25] LWL[24] LWL[23] LWL[22] LWL[21] LWL[20] LWL[19]
+ RWL[23] RWL[24] RWL[27] RWL[30] RWL[31] LWL[31] LWL[30] LWL[29] RWL[19] xa[2] xa[7]
+ xb[3] xb[2] xb[0] xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7219_n156# RWL[20] xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7483_n156#
+ xa[6] RWL[21] RWL[25] xa[3] xa[0] RWL[28] RWL[1] men xc xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7748_n156#
+ RWL[7] RWL[4] RWL[16] xa[5] RWL[9] RWL[29] RWL[22] xa[4] xb[1] RWL[15] RWL[26] xa[1]
+ RWL[12] vdd vss
Xxdec8_3v256x8m81_0 LWL[29] LWL[28] LWL[26] RWL[29] RWL[28] RWL[26] RWL[31] LWL[25]
+ LWL[31] LWL[30] LWL[24] LWL[27] xb[3] xa[4] xa[7] xa[1] xb[3] xb[3] xc xc xc xc
+ xb[3] xb[3] xa[3] xb[3] xa[0] xa[6] xa[7] RWL[27] xc xc xb[3] xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7219_n156#
+ xb[3] xa[3] xa[5] xa[2] RWL[24] xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7483_n156#
+ xa[0] RWL[30] xa[2] xa[6] xb[0] men xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7748_n156#
+ xa[4] xb[2] xa[1] xb[3] RWL[25] xb[1] xc xc vdd vss xa[5] xc xdec8_3v256x8m81
Xxdec8_3v256x8m81_1 LWL[5] LWL[4] LWL[2] RWL[5] RWL[4] RWL[2] RWL[7] LWL[1] LWL[7]
+ LWL[6] LWL[0] LWL[3] xb[0] xa[4] xa[7] xa[1] xb[0] xb[0] xc xc xc xc xb[0] xb[0]
+ xa[3] xb[0] xa[0] xa[6] xa[7] RWL[3] xc xc xb[0] xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7219_n156#
+ xb[0] xa[3] xa[5] xa[2] RWL[0] xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7483_n156#
+ xa[0] RWL[6] xa[2] xa[6] xb[0] men xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7748_n156#
+ xa[4] xb[2] xa[1] xb[3] RWL[1] xb[1] xc xc vdd vss xa[5] xc xdec8_3v256x8m81
Xxdec8_3v256x8m81_2 LWL[13] LWL[12] LWL[10] RWL[13] RWL[12] RWL[10] RWL[15] LWL[9]
+ LWL[15] LWL[14] LWL[8] LWL[11] xb[1] xa[4] xa[7] xa[1] xb[1] xb[1] xc xc xc xc xb[1]
+ xb[1] xa[3] xb[1] xa[0] xa[6] xa[7] RWL[11] xc xc xb[1] xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7219_n156#
+ xb[1] xa[3] xa[5] xa[2] RWL[8] xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7483_n156#
+ xa[0] RWL[14] xa[2] xa[6] xb[0] men xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7748_n156#
+ xa[4] xb[2] xa[1] xb[3] RWL[9] xb[1] xc xc vdd vss xa[5] xc xdec8_3v256x8m81
Xxdec8_3v256x8m81_3 LWL[21] LWL[20] LWL[18] RWL[21] RWL[20] RWL[18] RWL[23] LWL[17]
+ LWL[23] LWL[22] LWL[16] LWL[19] xb[2] xa[4] xa[7] xa[1] xb[2] xb[2] xc xc xc xc
+ xb[2] xb[2] xa[3] xb[2] xa[0] xa[6] xa[7] RWL[19] xc xc xb[2] xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7219_n156#
+ xb[2] xa[3] xa[5] xa[2] RWL[16] xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7483_n156#
+ xa[0] RWL[22] xa[2] xa[6] xb[0] men xdec8_3v256x8m81_3/xdec_3v256x8m81_7/m2_7748_n156#
+ xa[4] xb[2] xa[1] xb[3] RWL[17] xb[1] xc xc vdd vss xa[5] xc xdec8_3v256x8m81
.ends

.subckt pmos_5p043105913020100_3v256x8m81 D a_n28_n44# a_132_n44# w_n202_n86# S_uq0
+ S
X0 D a_n28_n44# S w_n202_n86# pfet_03v3 ad=1.5314p pd=6.41u as=2.5916p ps=12.66u w=5.89u l=0.28u
X1 S_uq0 a_132_n44# D w_n202_n86# pfet_03v3 ad=2.5916p pd=12.66u as=1.5314p ps=6.41u w=5.89u l=0.28u
.ends

.subckt pmos_1p2_02_R90_3v256x8m81 pmos_5p043105913020100_3v256x8m81_0/D w_n138_n63#
+ a_118_n33# pmos_5p043105913020100_3v256x8m81_0/S a_n41_n33# pmos_5p043105913020100_3v256x8m81_0/S_uq0
Xpmos_5p043105913020100_3v256x8m81_0 pmos_5p043105913020100_3v256x8m81_0/D a_n41_n33#
+ a_118_n33# w_n138_n63# pmos_5p043105913020100_3v256x8m81_0/S_uq0 pmos_5p043105913020100_3v256x8m81_0/S
+ pmos_5p043105913020100_3v256x8m81
.ends

.subckt nmos_5p04310591302099_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=2.0746p pd=10.31u as=2.0746p ps=10.31u w=4.715u l=0.28u
.ends

.subckt nmos_5p043105913020111_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=0.5412p pd=3.34u as=0.5412p ps=3.34u w=1.23u l=0.28u
.ends

.subckt pmoscap_R270_3v256x8m81 m3_770_16# a_n126_928# a_n140_236# m3_152_0# w_n226_n219#
X0 a_n140_236# a_n126_928# a_n140_236# w_n226_n219# pfet_03v3 ad=1.20555p pd=6.07u as=0 ps=0 w=2.565u l=2.505u
X1 a_n140_236# a_n126_928# a_n140_236# w_n226_n219# pfet_03v3 ad=0.6733p pd=3.09u as=0 ps=0 w=2.565u l=2.505u
.ends

.subckt nmos_1p2_02_R90_3v256x8m81 nmos_5p04310591302099_3v256x8m81_0/D a_n14_n33#
+ nmos_5p04310591302099_3v256x8m81_0/S VSUBS
Xnmos_5p04310591302099_3v256x8m81_0 nmos_5p04310591302099_3v256x8m81_0/D a_n14_n33#
+ nmos_5p04310591302099_3v256x8m81_0/S VSUBS nmos_5p04310591302099_3v256x8m81
.ends

.subckt pmoscap_L1_W2_R270_3v256x8m81 m3_307_0# m3_600_0# M2_M1$04_R270_3v256x8m81_0/VSUBS
+ a_597_236# m1_38_36# a_8_236#
X0 a_597_236# M2_M1$04_R270_3v256x8m81_0/VSUBS a_8_236# m1_38_36# pfet_03v3 ad=1.1286p pd=6.01u as=1.1286p ps=6.01u w=2.565u l=2.505u
.ends

.subckt nmos_5p043105913020102_3v256x8m81 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_03v3 ad=1.353p pd=7.03u as=1.353p ps=7.03u w=3.075u l=0.28u
.ends

.subckt nmos_1p2_01_R270_3v256x8m81 nmos_5p043105913020102_3v256x8m81_0/D a_n14_n33#
+ VSUBS nmos_5p043105913020102_3v256x8m81_0/S
Xnmos_5p043105913020102_3v256x8m81_0 nmos_5p043105913020102_3v256x8m81_0/D a_n14_n33#
+ nmos_5p043105913020102_3v256x8m81_0/S VSUBS nmos_5p043105913020102_3v256x8m81
.ends

.subckt pmos_1p2_01_R90_3v256x8m81 pmos_5p043105913020101_3v256x8m81_0/S w_n137_n63#
+ pmos_5p043105913020101_3v256x8m81_0/D a_n14_n33#
Xpmos_5p043105913020101_3v256x8m81_0 pmos_5p043105913020101_3v256x8m81_0/D a_n14_n33#
+ w_n137_n63# pmos_5p043105913020101_3v256x8m81_0/S pmos_5p043105913020101_3v256x8m81
.ends

.subckt xdec64_3v256x8m81 DRWL DLWL LWL[20] LWL[21] LWL[22] LWL[27] LWL[13] LWL[14]
+ LWL[16] LWL[3] LWL[2] LWL[1] LWL[0] LWL[8] LWL[9] LWL[7] LWL[30] RWL[31] RWL[30]
+ RWL[29] RWL[22] RWL[4] RWL[2] RWL[0] RWL[1] RWL[3] RWL[7] RWL[9] RWL[11] RWL[14]
+ RWL[15] RWL[16] RWL[17] RWL[18] RWL[19] RWL[20] xb[0] xb[1] xb[2] xb[3] xa[7] xa[6]
+ xa[5] xa[4] xa[0] men xa[3] xa[2] xa[1] xc[0] xc[1] RWL[21] LWL[25] LWL[28] LWL[26]
+ LWL[11] LWL[12] LWL[24] RWL[27] LWL[23] LWL[10] LWL[31] LWL[19] RWL[12] LWL[17]
+ RWL[28] RWL[25] RWL[10] LWL[29] RWL[5] RWL[26] LWL[5] LWL[6] RWL[13] LWL[18] RWL[24]
+ RWL[8] LWL[4] LWL[15] vdd vss RWL[23] RWL[6]
Xpmos_5p043105913020101_3v256x8m81_0 vdd pmos_5p043105913020101_3v256x8m81_1/D vdd
+ pmos_5p043105913020101_3v256x8m81_0/S pmos_5p043105913020101_3v256x8m81
Xpmos_5p043105913020101_3v256x8m81_1 pmos_5p043105913020101_3v256x8m81_1/D vss vdd
+ men pmos_5p043105913020101_3v256x8m81
Xxdec32_3v256x8m81_0 LWL[6] LWL[7] RWL[18] RWL[17] RWL[14] RWL[13] LWL[9] LWL[8] LWL[0]
+ LWL[1] LWL[2] LWL[3] LWL[4] LWL[5] RWL[11] RWL[10] RWL[8] RWL[5] RWL[3] RWL[0] RWL[2]
+ LWL[18] LWL[17] LWL[16] LWL[15] LWL[14] LWL[13] LWL[12] LWL[11] LWL[10] RWL[6] LWL[28]
+ LWL[27] LWL[26] LWL[25] LWL[24] LWL[23] LWL[22] LWL[21] LWL[20] LWL[19] RWL[23]
+ RWL[24] RWL[27] RWL[30] RWL[31] LWL[31] LWL[30] LWL[29] RWL[19] xa[2] xa[7] xb[3]
+ xb[2] xb[0] vdd RWL[20] vdd xa[6] RWL[21] RWL[25] xa[3] xa[0] RWL[28] RWL[1] men
+ xc[0] xc[1] RWL[7] RWL[4] RWL[16] xa[5] RWL[9] RWL[29] RWL[22] xa[4] xb[1] RWL[15]
+ RWL[26] xa[1] RWL[12] vdd vss xdec32_3v256x8m81
Xpmos_1p2_02_R90_3v256x8m81_0 DLWL vdd nmos_5p043105913020111_3v256x8m81_0/S vdd nmos_5p043105913020111_3v256x8m81_0/S
+ vdd pmos_1p2_02_R90_3v256x8m81
Xpmos_1p2_02_R90_3v256x8m81_1 DRWL vdd pmos_5p043105913020101_3v256x8m81_0/S vdd pmos_5p043105913020101_3v256x8m81_0/S
+ vdd pmos_1p2_02_R90_3v256x8m81
Xnmos_5p04310591302099_3v256x8m81_0 vss pmos_5p043105913020101_3v256x8m81_0/S DRWL
+ vss nmos_5p04310591302099_3v256x8m81
Xnmos_5p043105913020111_3v256x8m81_0 vss pmos_5p043105913020101_3v256x8m81_1/D nmos_5p043105913020111_3v256x8m81_0/S
+ vss nmos_5p043105913020111_3v256x8m81
Xnmos_5p043105913020111_3v256x8m81_1 vss pmos_5p043105913020101_3v256x8m81_1/D pmos_5p043105913020101_3v256x8m81_0/S
+ vss nmos_5p043105913020111_3v256x8m81
Xpmoscap_R270_3v256x8m81_0 RWL[16] vss vdd RWL[17] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_1 RWL[14] vss vdd RWL[15] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_2 RWL[12] vss vdd RWL[13] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_3 RWL[10] vss vdd RWL[11] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_4 RWL[8] vss vdd RWL[9] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_5 RWL[6] vss vdd RWL[7] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_6 RWL[4] vss vdd RWL[5] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_7 RWL[2] vss vdd RWL[3] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_8 RWL[0] vss vdd RWL[1] vdd pmoscap_R270_3v256x8m81
Xnmos_1p2_02_R90_3v256x8m81_0 vss nmos_5p043105913020111_3v256x8m81_0/S DLWL vss nmos_1p2_02_R90_3v256x8m81
Xpmoscap_R270_3v256x8m81_9 RWL[30] vss vdd RWL[31] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_30 LWL[20] vss vdd LWL[21] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_31 LWL[18] vss vdd LWL[19] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_20 LWL[8] vss vdd LWL[9] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_10 RWL[28] vss vdd RWL[29] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_21 LWL[6] vss vdd LWL[7] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_11 RWL[26] vss vdd RWL[27] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_22 LWL[4] vss vdd LWL[5] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_12 RWL[24] vss vdd RWL[25] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_23 LWL[2] vss vdd LWL[3] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_13 RWL[22] vss vdd RWL[23] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_24 LWL[0] vss vdd LWL[1] vdd pmoscap_R270_3v256x8m81
Xpmoscap_L1_W2_R270_3v256x8m81_0 DLWL vdd vss vdd vdd vdd pmoscap_L1_W2_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_25 LWL[30] vss vdd LWL[31] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_14 RWL[20] vss vdd RWL[21] vdd pmoscap_R270_3v256x8m81
Xpmoscap_L1_W2_R270_3v256x8m81_1 DRWL vdd vss vdd vdd vdd pmoscap_L1_W2_R270_3v256x8m81
Xnmos_1p2_01_R270_3v256x8m81_0 men vdd vss pmos_5p043105913020101_3v256x8m81_1/D nmos_1p2_01_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_26 LWL[28] vss vdd LWL[29] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_15 RWL[18] vss vdd RWL[19] vdd pmoscap_R270_3v256x8m81
Xpmos_1p2_01_R90_3v256x8m81_0 nmos_5p043105913020111_3v256x8m81_0/S vdd vdd pmos_5p043105913020101_3v256x8m81_1/D
+ pmos_1p2_01_R90_3v256x8m81
Xpmoscap_R270_3v256x8m81_27 LWL[26] vss vdd LWL[27] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_16 LWL[16] vss vdd LWL[17] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_28 LWL[24] vss vdd LWL[25] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_29 LWL[22] vss vdd LWL[23] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_17 LWL[14] vss vdd LWL[15] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_18 LWL[12] vss vdd LWL[13] vdd pmoscap_R270_3v256x8m81
Xpmoscap_R270_3v256x8m81_19 LWL[10] vss vdd LWL[11] vdd pmoscap_R270_3v256x8m81
.ends

.subckt gf180mcu_ocd_ip_sram__sram256x8m8wm1 A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0]
+ CEN CLK D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] GWEN Q[7] Q[6] Q[5] Q[4] Q[3] Q[2]
+ Q[1] Q[0] VDD VSS WEN[7] WEN[6] WEN[5] WEN[4] WEN[3] WEN[2] WEN[1] WEN[0]
Xlcol4_256_3v256x8m81_0 lcol4_256_3v256x8m81_0/WL[20] xdec64_3v256x8m81_0/LWL[20]
+ lcol4_256_3v256x8m81_0/WL[18] VSS VSS lcol4_256_3v256x8m81_0/WL[13] VSS VSS xdec64_3v256x8m81_0/LWL[9]
+ lcol4_256_3v256x8m81_0/WL[8] xdec64_3v256x8m81_0/LWL[7] lcol4_256_3v256x8m81_0/WL[6]
+ xdec64_3v256x8m81_0/LWL[5] xdec64_3v256x8m81_0/LWL[4] xdec64_3v256x8m81_0/LWL[3]
+ xdec64_3v256x8m81_0/LWL[2] xdec64_3v256x8m81_0/LWL[1] lcol4_256_3v256x8m81_0/WL[31]
+ lcol4_256_3v256x8m81_0/din[1] lcol4_256_3v256x8m81_0/din[3] lcol4_256_3v256x8m81_0/din[2]
+ lcol4_256_3v256x8m81_0/q[1] lcol4_256_3v256x8m81_0/q[2] lcol4_256_3v256x8m81_0/q[3]
+ lcol4_256_3v256x8m81_0/pcb[2] lcol4_256_3v256x8m81_0/pcb[3] lcol4_256_3v256x8m81_0/pcb[0]
+ lcol4_256_3v256x8m81_0/pcb[1] WEN[0] WEN[1] WEN[2] WEN[3] rcol4_256_3v256x8m81_0/GWE
+ Q[0] Q[1] control_3v256x8_3v256x8m81_0/IGWEN xdec64_3v256x8m81_0/LWL[6] xdec64_3v256x8m81_0/LWL[8]
+ xdec64_3v256x8m81_0/LWL[21] D[1] xdec64_3v256x8m81_0/LWL[22] VDD xdec64_3v256x8m81_0/LWL[23]
+ xdec64_3v256x8m81_0/LWL[24] xdec64_3v256x8m81_0/LWL[25] xdec64_3v256x8m81_0/LWL[26]
+ xdec64_3v256x8m81_0/LWL[27] D[3] xdec64_3v256x8m81_0/LWL[28] D[2] xdec64_3v256x8m81_0/LWL[29]
+ Q[3] Q[2] control_3v256x8_3v256x8m81_0/LYS[7] lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[1]
+ lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[2] rcol4_256_3v256x8m81_0/GWE
+ control_3v256x8_3v256x8m81_0/VDD_uq4 rcol4_256_3v256x8m81_0/GWE D[0] lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[4]
+ xdec64_3v256x8m81_0/men xdec64_3v256x8m81_0/LWL[10] lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[5]
+ xdec64_3v256x8m81_0/LWL[11] lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[6]
+ lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[7] xdec64_3v256x8m81_0/LWL[12]
+ rcol4_256_3v256x8m81_0/GWE VDD xdec64_3v256x8m81_0/LWL[30] xdec64_3v256x8m81_0/LWL[13]
+ VDD xdec64_3v256x8m81_0/LWL[14] xdec64_3v256x8m81_0/LWL[31] VDD xdec64_3v256x8m81_0/LWL[15]
+ VDD xdec64_3v256x8m81_0/LWL[16] VDD xdec64_3v256x8m81_0/LWL[17] VDD xdec64_3v256x8m81_0/LWL[18]
+ rcol4_256_3v256x8m81_0/GWE xdec64_3v256x8m81_0/LWL[0] VSS xdec64_3v256x8m81_0/LWL[19]
+ VDD VDD lcol4_256_3v256x8m81
Xrcol4_256_3v256x8m81_0 xdec64_3v256x8m81_0/RWL[30] rcol4_256_3v256x8m81_0/WL[20]
+ xdec64_3v256x8m81_0/RWL[28] xdec64_3v256x8m81_0/RWL[31] rcol4_256_3v256x8m81_0/WL[18]
+ xdec64_3v256x8m81_0/RWL[16] rcol4_256_3v256x8m81_0/WL[31] rcol4_256_3v256x8m81_0/WL[14]
+ rcol4_256_3v256x8m81_0/WL[16] xdec64_3v256x8m81_0/RWL[27] xdec64_3v256x8m81_0/RWL[20]
+ xdec64_3v256x8m81_0/RWL[29] rcol4_256_3v256x8m81_0/WL[12] rcol4_256_3v256x8m81_0/WL[8]
+ xdec64_3v256x8m81_0/RWL[5] rcol4_256_3v256x8m81_0/WL[10] rcol4_256_3v256x8m81_0/WL[13]
+ rcol4_256_3v256x8m81_0/WL[6] rcol4_256_3v256x8m81_0/tblhl rcol4_256_3v256x8m81_0/GWE
+ xdec64_3v256x8m81_0/RWL[11] rcol4_256_3v256x8m81_0/din[7] rcol4_256_3v256x8m81_0/q[5]
+ rcol4_256_3v256x8m81_0/q[6] rcol4_256_3v256x8m81_0/q[7] rcol4_256_3v256x8m81_0/din[5]
+ rcol4_256_3v256x8m81_0/din[6] rcol4_256_3v256x8m81_0/q[4] rcol4_256_3v256x8m81_0/pcb[6]
+ rcol4_256_3v256x8m81_0/pcb[7] rcol4_256_3v256x8m81_0/pcb[4] WEN[7] WEN[4] rcol4_256_3v256x8m81_0/pcb[5]
+ WEN[6] WEN[5] xdec64_3v256x8m81_0/RWL[17] rcol4_256_3v256x8m81_0/saout_R_m2_3v256x8m81_1/sa_3v256x8m81_0/pcb
+ xdec64_3v256x8m81_0/RWL[14] xdec64_3v256x8m81_0/RWL[13] control_3v256x8_3v256x8m81_0/RYS[1]
+ D[6] xdec64_3v256x8m81_0/men D[7] Q[6] xdec64_3v256x8m81_0/RWL[21] control_3v256x8_3v256x8m81_0/RYS[6]
+ xdec64_3v256x8m81_0/RWL[19] xdec64_3v256x8m81_0/RWL[15] control_3v256x8_3v256x8m81_0/RYS[7]
+ rcol4_256_3v256x8m81_0/saout_R_m2_3v256x8m81_1/sa_3v256x8m81_0/pcb VSS control_3v256x8_3v256x8m81_0/RYS[2]
+ xdec64_3v256x8m81_0/RWL[8] xdec64_3v256x8m81_0/RWL[22] xdec64_3v256x8m81_0/RWL[7]
+ xdec64_3v256x8m81_0/RWL[6] xdec64_3v256x8m81_0/RWL[1] xdec64_3v256x8m81_0/RWL[0]
+ control_3v256x8_3v256x8m81_0/RYS[0] xdec64_3v256x8m81_0/DRWL VDD xdec64_3v256x8m81_0/RWL[10]
+ VDD xdec64_3v256x8m81_0/RWL[9] xdec64_3v256x8m81_0/RWL[24] xdec64_3v256x8m81_0/RWL[23]
+ control_3v256x8_3v256x8m81_0/RYS[5] Q[7] Q[4] xdec64_3v256x8m81_0/RWL[2] control_3v256x8_3v256x8m81_0/RYS[4]
+ VDD VDD Q[5] D[5] xdec64_3v256x8m81_0/RWL[12] xdec64_3v256x8m81_0/RWL[26] VDD control_3v256x8_3v256x8m81_0/IGWEN
+ control_3v256x8_3v256x8m81_0/RYS[3] xdec64_3v256x8m81_0/RWL[25] VDD D[4] xdec64_3v256x8m81_0/RWL[4]
+ xdec64_3v256x8m81_0/RWL[3] xdec64_3v256x8m81_0/RWL[18] VDD VSS VDD rcol4_256_3v256x8m81
Xcontrol_3v256x8_3v256x8m81_0 VDD control_3v256x8_3v256x8m81_0/RYS[7] control_3v256x8_3v256x8m81_0/RYS[6]
+ control_3v256x8_3v256x8m81_0/RYS[5] control_3v256x8_3v256x8m81_0/RYS[4] control_3v256x8_3v256x8m81_0/RYS[3]
+ control_3v256x8_3v256x8m81_0/RYS[2] control_3v256x8_3v256x8m81_0/RYS[1] control_3v256x8_3v256x8m81_0/RYS[0]
+ VSS control_3v256x8_3v256x8m81_0/LYS[1] control_3v256x8_3v256x8m81_0/LYS[2] control_3v256x8_3v256x8m81_0/LYS[3]
+ control_3v256x8_3v256x8m81_0/LYS[6] control_3v256x8_3v256x8m81_0/LYS[5] control_3v256x8_3v256x8m81_0/LYS[4]
+ control_3v256x8_3v256x8m81_0/LYS[7] rcol4_256_3v256x8m81_0/tblhl control_3v256x8_3v256x8m81_0/IGWEN
+ xdec64_3v256x8m81_0/xb[3] xdec64_3v256x8m81_0/xb[2] xdec64_3v256x8m81_0/xb[0] xdec64_3v256x8m81_0/xa[7]
+ xdec64_3v256x8m81_0/xa[6] xdec64_3v256x8m81_0/xa[5] xdec64_3v256x8m81_0/xa[4] xdec64_3v256x8m81_0/xa[2]
+ A[0] xdec64_3v256x8m81_0/xb[1] control_3v256x8_3v256x8m81_0/xc[3] xdec64_3v256x8m81_0/xc[1]
+ control_3v256x8_3v256x8m81_0/xc[2] xdec64_3v256x8m81_0/xa[1] VSS A[7] CLK A[2] A[1]
+ A[6] A[3] A[4] A[5] VSS rcol4_256_3v256x8m81_0/GWE GWEN control_3v256x8_3v256x8m81_0/VSS_uq2
+ control_3v256x8_3v256x8m81_0/VSS_uq5 control_3v256x8_3v256x8m81_0/VDD_uq0 control_3v256x8_3v256x8m81_0/VDD_uq5
+ lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[1] lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[2]
+ xdec64_3v256x8m81_0/men control_3v256x8_3v256x8m81_0/VDD_uq4 lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[4]
+ xdec64_3v256x8m81_0/xa[3] lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[5]
+ lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[6] xdec64_3v256x8m81_0/xa[0]
+ lcol4_256_3v256x8m81_0/col_256a_3v256x8m81_0/ypass[7] CEN VDD VDD VDD control_3v256x8_3v256x8m81_0/xc[0]
+ VDD VDD VSS VDD VDD control_3v256x8_3v256x8m81
Xxdec64_3v256x8m81_0 xdec64_3v256x8m81_0/DRWL xdec64_3v256x8m81_0/DLWL xdec64_3v256x8m81_0/LWL[20]
+ xdec64_3v256x8m81_0/LWL[21] xdec64_3v256x8m81_0/LWL[22] xdec64_3v256x8m81_0/LWL[27]
+ xdec64_3v256x8m81_0/LWL[13] xdec64_3v256x8m81_0/LWL[14] xdec64_3v256x8m81_0/LWL[16]
+ xdec64_3v256x8m81_0/LWL[3] xdec64_3v256x8m81_0/LWL[2] xdec64_3v256x8m81_0/LWL[1]
+ xdec64_3v256x8m81_0/LWL[0] xdec64_3v256x8m81_0/LWL[8] xdec64_3v256x8m81_0/LWL[9]
+ xdec64_3v256x8m81_0/LWL[7] xdec64_3v256x8m81_0/LWL[30] xdec64_3v256x8m81_0/RWL[31]
+ xdec64_3v256x8m81_0/RWL[30] xdec64_3v256x8m81_0/RWL[29] xdec64_3v256x8m81_0/RWL[22]
+ xdec64_3v256x8m81_0/RWL[4] xdec64_3v256x8m81_0/RWL[2] xdec64_3v256x8m81_0/RWL[0]
+ xdec64_3v256x8m81_0/RWL[1] xdec64_3v256x8m81_0/RWL[3] xdec64_3v256x8m81_0/RWL[7]
+ xdec64_3v256x8m81_0/RWL[9] xdec64_3v256x8m81_0/RWL[11] xdec64_3v256x8m81_0/RWL[14]
+ xdec64_3v256x8m81_0/RWL[15] xdec64_3v256x8m81_0/RWL[16] xdec64_3v256x8m81_0/RWL[17]
+ xdec64_3v256x8m81_0/RWL[18] xdec64_3v256x8m81_0/RWL[19] xdec64_3v256x8m81_0/RWL[20]
+ xdec64_3v256x8m81_0/xb[0] xdec64_3v256x8m81_0/xb[1] xdec64_3v256x8m81_0/xb[2] xdec64_3v256x8m81_0/xb[3]
+ xdec64_3v256x8m81_0/xa[7] xdec64_3v256x8m81_0/xa[6] xdec64_3v256x8m81_0/xa[5] xdec64_3v256x8m81_0/xa[4]
+ xdec64_3v256x8m81_0/xa[0] xdec64_3v256x8m81_0/men xdec64_3v256x8m81_0/xa[3] xdec64_3v256x8m81_0/xa[2]
+ xdec64_3v256x8m81_0/xa[1] VDD xdec64_3v256x8m81_0/xc[1] xdec64_3v256x8m81_0/RWL[21]
+ xdec64_3v256x8m81_0/LWL[25] xdec64_3v256x8m81_0/LWL[28] xdec64_3v256x8m81_0/LWL[26]
+ xdec64_3v256x8m81_0/LWL[11] xdec64_3v256x8m81_0/LWL[12] xdec64_3v256x8m81_0/LWL[24]
+ xdec64_3v256x8m81_0/RWL[27] xdec64_3v256x8m81_0/LWL[23] xdec64_3v256x8m81_0/LWL[10]
+ xdec64_3v256x8m81_0/LWL[31] xdec64_3v256x8m81_0/LWL[19] xdec64_3v256x8m81_0/RWL[12]
+ xdec64_3v256x8m81_0/LWL[17] xdec64_3v256x8m81_0/RWL[28] xdec64_3v256x8m81_0/RWL[25]
+ xdec64_3v256x8m81_0/RWL[10] xdec64_3v256x8m81_0/LWL[29] xdec64_3v256x8m81_0/RWL[5]
+ xdec64_3v256x8m81_0/RWL[26] xdec64_3v256x8m81_0/LWL[5] xdec64_3v256x8m81_0/LWL[6]
+ xdec64_3v256x8m81_0/RWL[13] xdec64_3v256x8m81_0/LWL[18] xdec64_3v256x8m81_0/RWL[24]
+ xdec64_3v256x8m81_0/RWL[8] xdec64_3v256x8m81_0/LWL[4] xdec64_3v256x8m81_0/LWL[15]
+ VDD VSS xdec64_3v256x8m81_0/RWL[23] xdec64_3v256x8m81_0/RWL[6] xdec64_3v256x8m81
.ends

