magic
tech gf180mcuD
magscale 1 10
timestamp 1763578215
<< metal2 >>
rect -4 2229 151 13188
rect 346 2891 503 11480
rect 707 2229 863 13180
use M2_M14310591302097_512x8m81  M2_M14310591302097_512x8m81_0
timestamp 1763564386
transform 1 0 784 0 1 2560
box -70 -330 70 330
use M2_M14310591302097_512x8m81  M2_M14310591302097_512x8m81_1
timestamp 1763564386
transform 1 0 72 0 1 2560
box -70 -330 70 330
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_0
timestamp 1763564386
transform 1 0 424 0 1 5145
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_1
timestamp 1763564386
transform 1 0 786 0 1 3898
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_2
timestamp 1763564386
transform 1 0 74 0 1 4687
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_3
timestamp 1763564386
transform 1 0 786 0 1 4687
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_4
timestamp 1763564386
transform 1 0 424 0 1 5739
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_5
timestamp 1763564386
transform 1 0 786 0 1 6138
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_6
timestamp 1763564386
transform 1 0 74 0 1 6138
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_7
timestamp 1763564386
transform 1 0 74 0 1 3898
box -70 -113 70 113
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_0
timestamp 1763564386
transform 1 0 74 0 1 6968
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_1
timestamp 1763564386
transform 1 0 74 0 1 9451
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_2
timestamp 1763564386
transform 1 0 786 0 1 9451
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_3
timestamp 1763564386
transform 1 0 74 0 1 8970
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_4
timestamp 1763564386
transform 1 0 786 0 1 8970
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_5
timestamp 1763564386
transform 1 0 74 0 1 12935
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_6
timestamp 1763564386
transform 1 0 786 0 1 12935
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_7
timestamp 1763564386
transform 1 0 74 0 1 12454
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_8
timestamp 1763564386
transform 1 0 786 0 1 12454
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_9
timestamp 1763564386
transform 1 0 74 0 1 11975
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_10
timestamp 1763564386
transform 1 0 786 0 1 11975
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_11
timestamp 1763564386
transform 1 0 786 0 1 6968
box -70 -200 70 200
use M3_M24310591302099_512x8m81  M3_M24310591302099_512x8m81_0
timestamp 1763564386
transform 1 0 424 0 1 10800
box -70 -634 70 634
use M3_M243105913020100_512x8m81  M3_M243105913020100_512x8m81_0
timestamp 1763564386
transform 1 0 424 0 1 7792
box -70 -417 70 417
use M3_M243105913020101_512x8m81  M3_M243105913020101_512x8m81_0
timestamp 1763564386
transform 1 0 424 0 1 3233
box -70 -330 70 330
<< end >>
