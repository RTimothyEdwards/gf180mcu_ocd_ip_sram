magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal3 >>
rect -357 441 342 1701
use M3_M24310591302042_512x8m81  M3_M24310591302042_512x8m81_0
timestamp 1763564386
transform 1 0 -8 0 1 788
box -330 -330 330 330
<< properties >>
string path -0.055 3.150 -0.055 12.150 
<< end >>
