magic
tech gf180mcuD
magscale 1 10
timestamp 1765833244
<< nwell >>
rect -174 -86 230 1144
<< pmos >>
rect 0 0 56 1058
<< pdiff >>
rect -88 1045 0 1058
rect -88 13 -75 1045
rect -29 13 0 1045
rect -88 0 0 13
rect 56 1045 144 1058
rect 56 13 85 1045
rect 131 13 144 1045
rect 56 0 144 13
<< pdiffc >>
rect -75 13 -29 1045
rect 85 13 131 1045
<< polysilicon >>
rect 0 1058 56 1102
rect 0 -44 56 0
<< metal1 >>
rect -75 1045 -29 1058
rect -75 0 -29 13
rect 85 1045 131 1058
rect 85 0 131 13
<< labels >>
flabel pdiffc -40 529 -40 529 0 FreeSans 186 0 0 0 S
flabel pdiffc 96 529 96 529 0 FreeSans 186 0 0 0 D
<< end >>
