magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< psubdiff >>
rect -2655 23 2635 56
rect -2655 -23 -2624 23
rect 2604 -23 2635 23
rect -2655 -56 2635 -23
<< psubdiffcont >>
rect -2624 -23 2604 23
<< metal1 >>
rect -2641 23 2621 42
rect -2641 -23 -2624 23
rect 2604 -23 2621 23
rect -2641 -42 2621 -23
<< end >>
