magic
tech gf180mcuD
magscale 1 10
timestamp 1764700137
<< nwell >>
rect 91 512 511 797
<< pwell >>
rect 91 55 511 512
<< psubdiff >>
rect 238 296 362 319
rect 238 150 277 296
rect 323 150 362 296
rect 238 55 362 150
<< nsubdiff >>
rect 138 758 462 773
rect 138 706 177 758
rect 423 706 462 758
rect 138 643 462 706
<< psubdiffcont >>
rect 277 150 323 296
<< nsubdiffcont >>
rect 177 706 423 758
<< polysilicon >>
rect 117 533 482 570
rect 117 487 177 533
rect 423 487 482 533
rect 117 450 482 487
rect 117 250 176 450
rect 91 178 176 250
rect 424 250 482 450
rect 424 178 511 250
<< polycontact >>
rect 177 487 423 533
<< metal1 >>
rect 91 758 511 760
rect 91 706 114 758
rect 166 706 177 758
rect 423 706 511 758
rect 91 704 511 706
rect 228 644 372 646
rect 228 592 274 644
rect 326 592 372 644
rect 228 582 372 592
rect 118 536 482 582
rect 118 533 274 536
rect 326 533 482 536
rect 118 487 177 533
rect 423 487 482 533
rect 118 484 274 487
rect 326 484 482 487
rect 118 438 482 484
rect 228 428 372 438
rect 228 376 274 428
rect 326 376 372 428
rect 228 374 372 376
rect 91 296 511 321
rect 91 199 277 296
rect 218 150 277 199
rect 323 287 511 296
rect 323 235 434 287
rect 486 235 511 287
rect 323 199 511 235
rect 323 150 382 199
rect 218 89 382 150
<< via1 >>
rect 114 706 166 758
rect 274 592 326 644
rect 274 533 326 536
rect 274 487 326 533
rect 274 484 326 487
rect 274 376 326 428
rect 434 235 486 287
<< metal2 >>
rect 103 758 194 772
rect 103 706 114 758
rect 166 706 194 758
rect 103 55 194 706
rect 250 374 272 646
rect 328 374 350 646
rect 406 287 499 772
rect 406 235 434 287
rect 486 235 499 287
rect 406 55 499 235
<< via2 >>
rect 272 644 328 646
rect 272 592 274 644
rect 274 592 326 644
rect 326 592 328 644
rect 272 536 328 592
rect 272 484 274 536
rect 274 484 326 536
rect 326 484 328 536
rect 272 428 328 484
rect 272 376 274 428
rect 274 376 326 428
rect 326 376 328 428
rect 272 374 328 376
<< metal3 >>
rect 91 646 511 690
rect 91 374 272 646
rect 328 374 511 646
rect 91 330 511 374
rect 91 56 511 196
use M2_M14310591302020_3v256x8m81  M2_M14310591302020_3v256x8m81_0
timestamp 1764700137
transform 1 0 300 0 1 126
box -35 -56 35 55
use M3_M24310591302021_3v256x8m81  M3_M24310591302021_3v256x8m81_0
timestamp 1764700137
transform 1 0 300 0 1 126
box -35 -35 35 35
<< properties >>
string FIXED_BBOX -68 -68 668 968
string MASKHINTS_SRAMDEF 91 89 511 797
<< end >>
