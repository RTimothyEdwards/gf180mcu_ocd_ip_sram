magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< error_s >>
rect 1245 2672 1359 4262
<< nwell >>
rect 2849 7017 3760 7028
rect 2644 6920 3760 7017
rect 2644 6563 4661 6920
rect 2644 6554 3760 6563
rect 2650 5234 2999 5247
rect 2507 2629 2999 5234
rect 3728 3278 3877 5233
rect 3368 3262 3877 3278
rect 4176 3263 4953 5302
rect 3802 557 3850 1390
<< pmos >>
rect 3035 6653 3091 6813
rect 3195 6653 3251 6813
rect 3360 6653 3416 6813
rect 3497 6653 3553 6813
<< pdiff >>
rect 2944 6799 3035 6813
rect 2944 6678 2958 6799
rect 3004 6678 3035 6799
rect 2944 6653 3035 6678
rect 3091 6653 3195 6813
rect 3251 6799 3360 6813
rect 3251 6678 3280 6799
rect 3326 6678 3360 6799
rect 3251 6653 3360 6678
rect 3416 6653 3497 6813
rect 3553 6799 3665 6813
rect 3553 6678 3595 6799
rect 3642 6678 3665 6799
rect 3553 6653 3665 6678
<< pdiffc >>
rect 2958 6678 3004 6799
rect 3280 6678 3326 6799
rect 3595 6678 3642 6799
<< nsubdiff >>
rect 2609 5019 2807 5131
<< polysilicon >>
rect 3420 7237 3479 7324
rect 3035 6813 3091 7139
rect 3195 7126 3251 7139
rect 3390 7126 3449 7207
rect 3195 7051 3449 7126
rect 3195 6813 3251 7051
rect 3360 7044 3449 7051
rect 3360 6813 3416 7044
rect 3556 6976 3692 7035
rect 3497 6934 3692 6976
rect 3497 6813 3553 6934
rect 4151 6918 4207 7143
rect 4073 6864 4289 6918
rect 4073 6812 4129 6864
rect 4233 6812 4289 6864
rect 3035 6602 3091 6653
rect 3195 6602 3251 6653
rect 3360 6602 3416 6653
rect 3497 6602 3553 6653
rect 4073 6550 4129 6627
rect 4233 6550 4289 6628
<< metal1 >>
rect 2950 7920 3032 7975
rect 2950 7168 3031 7920
rect 3107 7106 3188 7301
rect 3264 7168 3345 7979
rect 4223 7920 4305 8003
rect 4223 7562 4304 7920
rect 3107 7023 3345 7106
rect 4076 7084 4123 7254
rect 4223 7221 4305 7562
rect 2950 6799 3031 6895
rect 2950 6678 2958 6799
rect 3004 6678 3031 6799
rect 2950 6659 3031 6678
rect 3264 6799 3345 7023
rect 3562 6955 3675 7026
rect 4076 6990 5013 7084
rect 3264 6678 3280 6799
rect 3326 6678 3345 6799
rect 3264 6603 3345 6678
rect 3577 6799 4041 6895
rect 3577 6678 3595 6799
rect 3642 6678 4041 6799
rect 4157 6731 4204 6990
rect 3577 6663 4041 6678
rect 4322 6668 4581 6895
rect 3577 6659 3658 6663
rect 3264 6519 4279 6603
rect 2806 5116 2893 5117
rect 2538 5033 2893 5116
rect 3213 2597 3304 2979
<< metal2 >>
rect 457 7739 548 7833
rect 706 7739 797 7833
rect 1710 7739 1801 7833
rect 1963 7739 2054 7833
rect 3402 7357 3493 7451
rect 2809 7014 3675 7108
rect 3773 6510 3864 6603
rect 3773 3831 3863 6510
rect 3413 3738 3863 3831
rect 3413 2571 3503 3738
rect 3573 2441 3663 3614
rect 4397 2314 4487 2979
rect 4757 2173 4847 3614
rect 4929 2981 5020 6981
rect 3612 148 3702 242
rect 4795 148 4886 242
<< metal3 >>
rect -202 7013 5166 7679
rect -202 6435 5166 6934
rect -202 5705 5166 6342
rect -202 3563 5166 5469
rect 289 1563 5166 2041
rect 289 754 5166 1390
rect 289 0 5166 634
use M1_NACTIVE4310591302028_512x8m81  M1_NACTIVE4310591302028_512x8m81_0
timestamp 1763476864
transform 1 0 2793 0 1 6776
box -36 -95 36 95
use M1_NACTIVE4310591302028_512x8m81  M1_NACTIVE4310591302028_512x8m81_1
timestamp 1763476864
transform 1 0 4537 0 1 6776
box -36 -95 36 95
use M1_PACTIVE_02_512x8m81  M1_PACTIVE_02_512x8m81_0
timestamp 1763476864
transform 1 0 3836 0 1 7963
box -1382 -56 1382 56
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_0
timestamp 1763476864
transform 1 0 2324 0 1 2488
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_1
timestamp 1763476864
transform 1 0 1065 0 1 2631
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_2
timestamp 1763476864
transform 1 0 1443 0 1 2488
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_3
timestamp 1763476864
transform 1 0 2163 0 1 2205
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_4
timestamp 1763476864
transform 1 0 345 0 1 2345
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_5
timestamp 1763476864
transform 1 0 868 0 1 2205
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_6
timestamp 1763476864
transform 1 0 179 0 1 2631
box -67 -48 67 47
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_7
timestamp 1763476864
transform 1 0 1605 0 1 2345
box -67 -48 67 47
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_0
timestamp 1763476864
transform 0 -1 2969 1 0 7055
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_1
timestamp 1763476864
transform 0 -1 3619 1 0 6971
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_2
timestamp 1763476864
transform 1 0 3449 0 1 7262
box -36 -126 60 122
use M1_POLY24310591302030_512x8m81  M1_POLY24310591302030_512x8m81_0
timestamp 1763476864
transform 1 0 4189 0 1 6586
box -95 -36 95 36
use M2_M1$$34864172_512x8m81  M2_M1$$34864172_512x8m81_0
timestamp 1763476864
transform 1 0 3818 0 1 6556
box -119 -46 119 46
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1763476864
transform 1 0 4975 0 1 6985
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_1
timestamp 1763476864
transform 1 0 2986 0 1 6763
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_2
timestamp 1763476864
transform 1 0 4536 0 1 6773
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_3
timestamp 1763476864
transform 1 0 2793 0 1 6763
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_4
timestamp 1763476864
transform 1 0 3448 0 1 7328
box -43 -122 43 122
use M2_M1$$43375660_R90_512x8m81  M2_M1$$43375660_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 3819 1 0 6722
box -46 -119 46 119
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_0
timestamp 1763476864
transform 1 0 2986 0 1 7403
box -44 -198 44 198
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_1
timestamp 1763476864
transform 1 0 3294 0 1 7403
box -44 -198 44 198
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_2
timestamp 1763476864
transform 1 0 4263 0 1 7363
box -44 -198 44 198
use M2_M1$$46894124_512x8m81  M2_M1$$46894124_512x8m81_0
timestamp 1763476864
transform 1 0 3618 0 1 2488
box -44 -46 45 46
use M2_M1$$46894124_512x8m81  M2_M1$$46894124_512x8m81_1
timestamp 1763476864
transform 1 0 4442 0 1 2347
box -44 -46 45 46
use M2_M1$$46894124_512x8m81  M2_M1$$46894124_512x8m81_2
timestamp 1763476864
transform 1 0 4802 0 1 2205
box -44 -46 45 46
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_0
timestamp 1763476864
transform 1 0 2963 0 1 7053
box -63 -34 63 34
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_1
timestamp 1763476864
transform 1 0 3612 0 1 7053
box -63 -34 63 34
use M3_M2$$43368492_R90_512x8m81  M3_M2$$43368492_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 3819 1 0 6722
box -46 -119 46 119
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_0
timestamp 1763476864
transform 1 0 2986 0 1 6687
box -45 -198 45 198
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_1
timestamp 1763476864
transform 1 0 4536 0 1 6696
box -45 -198 45 198
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_2
timestamp 1763476864
transform 1 0 2986 0 1 7403
box -45 -198 45 198
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_3
timestamp 1763476864
transform 1 0 3294 0 1 7403
box -45 -198 45 198
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_4
timestamp 1763476864
transform 1 0 2793 0 1 6687
box -45 -198 45 198
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_5
timestamp 1763476864
transform 1 0 4263 0 1 7363
box -45 -198 45 198
use nmos_1p2$$46563372_512x8m81  nmos_1p2$$46563372_512x8m81_0
timestamp 1763476864
transform 1 0 4165 0 1 7165
box -102 -44 130 133
use nmos_5p04310591302040_512x8m81  nmos_5p04310591302040_512x8m81_0
timestamp 1763476864
transform 1 0 3035 0 1 7168
box -88 -44 144 171
use nmos_5p04310591302040_512x8m81  nmos_5p04310591302040_512x8m81_1
timestamp 1763476864
transform 1 0 3195 0 1 7168
box -88 -44 144 171
use pmos_5p04310591302069_512x8m81  pmos_5p04310591302069_512x8m81_0
timestamp 1763476864
transform 1 0 4101 0 1 6663
box -202 -86 362 192
use xpredec0_bot_512x8m81  xpredec0_bot_512x8m81_0
timestamp 1763476864
transform 1 0 3796 0 1 442
box -74 -442 1276 5901
use xpredec0_bot_512x8m81  xpredec0_bot_512x8m81_1
timestamp 1763476864
transform 1 0 2613 0 1 442
box -74 -442 1276 5901
use xpredec0_xa_512x8m81  xpredec0_xa_512x8m81_0
timestamp 1763476864
transform -1 0 2817 0 1 23
box 107 -24 1143 7982
use xpredec0_xa_512x8m81  xpredec0_xa_512x8m81_1
timestamp 1763476864
transform -1 0 1537 0 1 23
box 107 -24 1143 7982
use xpredec0_xa_512x8m81  xpredec0_xa_512x8m81_2
timestamp 1763476864
transform 1 0 947 0 1 23
box 107 -24 1143 7982
use xpredec0_xa_512x8m81  xpredec0_xa_512x8m81_3
timestamp 1763476864
transform 1 0 -333 0 1 23
box 107 -24 1143 7982
<< labels >>
rlabel metal3 s 5068 6655 5068 6655 4 vdd
port 1 nsew
rlabel metal3 s 5068 7318 5068 7318 4 vss
port 2 nsew
rlabel metal3 s 5068 4495 5068 4495 4 vdd
port 1 nsew
rlabel metal3 s 5068 289 5068 289 4 vss
port 2 nsew
rlabel metal3 s 5068 1061 5068 1061 4 vdd
port 1 nsew
rlabel metal3 s 5068 1785 5068 1785 4 vss
port 2 nsew
rlabel metal3 s 5068 6010 5068 6010 4 vss
port 2 nsew
rlabel metal2 s 4837 195 4837 195 4 A[0]
port 3 nsew
rlabel metal2 s 2854 7065 2854 7065 4 men
port 4 nsew
rlabel metal2 s 2006 7786 2006 7786 4 x[0]
port 5 nsew
rlabel metal2 s 1752 7786 1752 7786 4 x[1]
port 6 nsew
rlabel metal2 s 751 7786 751 7786 4 x[2]
port 7 nsew
rlabel metal2 s 502 7786 502 7786 4 x[3]
port 8 nsew
rlabel metal2 s 3654 195 3654 195 4 A[1]
port 9 nsew
rlabel metal2 s 3448 7401 3448 7401 4 clk
port 10 nsew
<< end >>
