magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal1 >>
rect -44 407 44 427
rect -44 -407 -26 407
rect 26 -407 44 407
rect -44 -427 44 -407
<< via1 >>
rect -26 -407 26 407
<< metal2 >>
rect -44 407 44 427
rect -44 -407 -26 407
rect 26 -407 44 407
rect -44 -427 44 -407
<< end >>
