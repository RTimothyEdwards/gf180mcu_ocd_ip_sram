magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal2 >>
rect -119 400 119 427
rect -119 -400 -93 400
rect 93 -400 119 400
rect -119 -427 119 -400
<< via2 >>
rect -93 -400 93 400
<< metal3 >>
rect -119 400 119 427
rect -119 -400 -93 400
rect 93 -400 119 400
rect -119 -427 119 -400
<< end >>
