magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect -29 -2598 695 -2070
rect -100 -2930 774 -2598
rect -29 -3360 695 -2930
<< nmos >>
rect 145 -7127 201 -5962
rect 305 -7127 361 -5962
rect 465 -7127 521 -5962
<< ndiff >>
rect 54 -5975 145 -5962
rect 54 -7102 70 -5975
rect 116 -7102 145 -5975
rect 54 -7127 145 -7102
rect 201 -7127 305 -5962
rect 361 -7127 465 -5962
rect 521 -5975 618 -5962
rect 521 -7102 550 -5975
rect 597 -7102 618 -5975
rect 521 -7127 618 -7102
<< ndiffc >>
rect 70 -7102 116 -5975
rect 550 -7102 597 -5975
<< psubdiff >>
rect 0 137 674 171
rect 0 91 141 137
rect 519 91 674 137
rect 0 56 674 91
rect 0 -7313 674 -7279
rect 0 -7359 141 -7313
rect 519 -7359 674 -7313
rect 0 -7394 674 -7359
<< nsubdiff >>
rect 0 -2747 674 -2715
rect 0 -2793 133 -2747
rect 401 -2793 674 -2747
rect 0 -2827 674 -2793
<< psubdiffcont >>
rect 141 91 519 137
rect 141 -7359 519 -7313
<< nsubdiffcont >>
rect 133 -2793 401 -2747
<< polysilicon >>
rect 145 -780 201 -558
rect 305 -780 361 -558
rect 465 -780 521 -558
rect 145 -876 521 -780
rect 145 -884 201 -876
rect 305 -884 361 -876
rect 465 -884 521 -876
rect 145 -2558 201 -2026
rect 305 -2558 361 -2026
rect 465 -2558 521 -2026
rect 137 -2653 535 -2558
rect 145 -5962 201 -4458
rect 305 -5962 361 -4458
rect 465 -5962 521 -4458
rect 145 -7178 201 -7127
rect 305 -7178 361 -7127
rect 465 -7178 521 -7127
<< metal1 >>
rect 0 137 674 165
rect 0 91 141 137
rect 519 91 674 137
rect 0 -38 674 91
rect 60 -39 142 -38
rect 60 -175 141 -39
rect 374 -175 455 -38
rect 217 -784 298 -465
rect 531 -784 611 -462
rect 217 -867 611 -784
rect 217 -968 298 -867
rect 531 -968 611 -867
rect 66 -2060 124 -1920
rect 385 -2061 443 -1921
rect 139 -2647 611 -2564
rect 0 -2747 455 -2729
rect 0 -2793 133 -2747
rect 401 -2793 455 -2747
rect 0 -2812 455 -2793
rect 60 -3024 142 -2812
rect 374 -3025 455 -2812
rect 531 -3496 611 -2647
rect -40 -4571 714 -4506
rect -40 -4712 714 -4648
rect -40 -4853 714 -4789
rect -40 -4994 714 -4930
rect -40 -5135 714 -5071
rect -40 -5277 714 -5212
rect 60 -5460 141 -5387
rect 60 -5975 142 -5460
rect 60 -7102 70 -5975
rect 116 -7102 142 -5975
rect 60 -7183 142 -7102
rect 531 -5975 612 -5387
rect 531 -7102 550 -5975
rect 597 -6547 612 -5975
rect 597 -7102 611 -6547
rect 531 -7121 611 -7102
rect 56 -7184 146 -7183
rect 5 -7313 674 -7184
rect 5 -7359 141 -7313
rect 519 -7359 674 -7313
rect 5 -7387 674 -7359
<< metal2 >>
rect 147 -499 301 228
rect 213 -4414 616 -4168
rect 527 -5591 616 -4414
<< metal3 >>
rect -36 -436 774 228
rect -40 -3887 774 -1981
rect 0 -5886 674 -5409
rect -46 -7451 774 -6815
use M1_POLY24310591302060_512x8m81  M1_POLY24310591302060_512x8m81_0
timestamp 1763476864
transform 1 0 343 0 1 -2604
box -128 -36 128 36
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1763476864
transform 1 0 571 0 1 -4291
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_1
timestamp 1763476864
transform 1 0 258 0 1 -4291
box -43 -122 43 122
use M2_M1$$43376684_512x8m81  M2_M1$$43376684_512x8m81_0
timestamp 1763476864
transform 1 0 571 0 1 -5966
box -44 -579 44 579
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_0
timestamp 1763476864
transform 1 0 420 0 1 -130
box -44 -275 44 275
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_0
timestamp 1763476864
transform 1 0 93 0 1 -2218
box -44 -198 44 198
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_1
timestamp 1763476864
transform 1 0 415 0 1 -2218
box -44 -198 44 198
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_2
timestamp 1763476864
transform 1 0 256 0 1 -299
box -44 -198 44 198
use M2_M1$$47327276_512x8m81  M2_M1$$47327276_512x8m81_0
timestamp 1763476864
transform 1 0 93 0 1 -6420
box -45 -961 45 961
use M2_M1$$47515692_512x8m81  M2_M1$$47515692_512x8m81_0
timestamp 1763476864
transform 1 0 93 0 1 -3306
box -44 -504 44 504
use M2_M1$$47515692_512x8m81  M2_M1$$47515692_512x8m81_1
timestamp 1763476864
transform 1 0 412 0 1 -3306
box -44 -504 44 504
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_0
timestamp 1763476864
transform 1 0 93 0 1 -2218
box -45 -198 45 198
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_1
timestamp 1763476864
transform 1 0 415 0 1 -2218
box -45 -198 45 198
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_2
timestamp 1763476864
transform 1 0 93 0 1 -5658
box -45 -198 45 198
use M3_M2$$47332396_512x8m81  M3_M2$$47332396_512x8m81_0
timestamp 1763476864
transform 1 0 93 0 1 -3306
box -45 -504 45 504
use M3_M2$$47332396_512x8m81  M3_M2$$47332396_512x8m81_1
timestamp 1763476864
transform 1 0 412 0 1 -3306
box -45 -504 45 504
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_0
timestamp 1763476864
transform 1 0 93 0 1 -7106
box -45 -275 45 275
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_1
timestamp 1763476864
transform 1 0 420 0 1 -130
box -45 -275 45 275
use nmos_1p2$$47514668_512x8m81  nmos_1p2$$47514668_512x8m81_0
timestamp 1763476864
transform 1 0 159 0 -1 -95
box -102 -44 130 467
use nmos_1p2$$47514668_512x8m81  nmos_1p2$$47514668_512x8m81_1
timestamp 1763476864
transform 1 0 319 0 -1 -95
box -102 -44 130 467
use nmos_1p2$$47514668_512x8m81  nmos_1p2$$47514668_512x8m81_2
timestamp 1763476864
transform 1 0 479 0 -1 -95
box -102 -44 130 467
use pmos_1p2$$47512620_512x8m81  pmos_1p2$$47512620_512x8m81_0
timestamp 1763476864
transform 1 0 479 0 1 -4419
box -188 -86 216 1059
use pmos_1p2$$47512620_512x8m81  pmos_1p2$$47512620_512x8m81_1
timestamp 1763476864
transform 1 0 319 0 1 -4419
box -188 -86 216 1059
use pmos_1p2$$47512620_512x8m81  pmos_1p2$$47512620_512x8m81_2
timestamp 1763476864
transform 1 0 159 0 1 -4419
box -188 -86 216 1059
use pmos_1p2$$47513644_512x8m81  pmos_1p2$$47513644_512x8m81_0
timestamp 1763476864
transform 1 0 319 0 -1 -926
box -188 -86 216 1144
use pmos_1p2$$47513644_512x8m81  pmos_1p2$$47513644_512x8m81_1
timestamp 1763476864
transform 1 0 479 0 -1 -926
box -188 -86 216 1144
use pmos_1p2$$47513644_512x8m81  pmos_1p2$$47513644_512x8m81_2
timestamp 1763476864
transform 1 0 159 0 -1 -926
box -188 -86 216 1144
<< end >>
