magic
tech gf180mcuD
magscale 1 10
timestamp 1764700137
use 018SRAM_cell1_3v256x8m81  018SRAM_cell1_3v256x8m81_0
timestamp 1764700137
transform 1 0 0 0 -1 900
box 30 89 570 797
use 018SRAM_cell1_3v256x8m81  018SRAM_cell1_3v256x8m81_1
timestamp 1764700137
transform 1 0 0 0 1 648
box 30 89 570 797
<< end >>
