magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal1 >>
rect -63 91 63 99
rect -63 -91 -54 91
rect 54 -91 63 91
rect -63 -99 63 -91
<< via1 >>
rect -54 -91 54 91
<< metal2 >>
rect -63 91 63 99
rect -63 -91 -54 91
rect 54 -91 63 91
rect -63 -99 63 -91
<< end >>
