magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
use 018SRAM_cell1_512x8m81  018SRAM_cell1_512x8m81_0
timestamp 1763765945
transform 1 0 0 0 -1 900
box 62 89 538 797
use 018SRAM_cell1_512x8m81  018SRAM_cell1_512x8m81_1
timestamp 1763765945
transform 1 0 0 0 1 648
box 62 89 538 797
<< end >>
