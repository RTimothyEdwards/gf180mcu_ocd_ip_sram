magic
tech gf180mcuD
magscale 1 10
timestamp 1764700137
<< nwell >>
rect 283 723 397 948
<< polysilicon >>
rect 533 3876 589 4647
rect 893 3876 949 4647
<< metal1 >>
rect 226 5369 529 5472
rect 227 4674 529 5369
rect 605 4612 686 4717
rect 605 4528 901 4612
rect 245 2573 529 4466
rect 605 3740 686 4528
rect 965 3767 1045 4717
rect -9 2436 1367 2501
rect -9 2295 1367 2360
rect -9 2154 1367 2219
rect -9 2013 1367 2077
rect -9 1871 1367 1936
rect -9 1730 1367 1795
<< metal2 >>
rect 294 4921 529 5472
rect 294 951 385 4617
rect 800 989 890 2657
rect 1144 1130 1233 2839
rect 800 896 1233 989
<< metal3 >>
rect 0 4882 1313 5518
rect 0 3120 1330 4645
rect 4 2821 1232 2914
rect 10 2563 1232 2657
use alatch_3v256x8m81  alatch_3v256x8m81_0
timestamp 1764700137
transform 1 0 49 0 1 -442
box -63 409 1197 2033
use M1_NWELL14_3v256x8m81  M1_NWELL14_3v256x8m81_0
timestamp 1763766357
transform 1 0 233 0 1 3542
box -154 -1016 154 1016
use M1_POLY2$$46559276_3v256x8m81  M1_POLY2$$46559276_3v256x8m81_0
timestamp 1763766357
transform 1 0 805 0 1 4570
box -123 -48 123 48
use M1_POLY2$$46559276_3v256x8m81  M1_POLY2$$46559276_3v256x8m81_1
timestamp 1763766357
transform 1 0 448 0 1 4570
box -123 -48 123 48
use M1_PSUB$$47818796_3v256x8m81  M1_PSUB$$47818796_3v256x8m81_0
timestamp 1763766357
transform 1 0 276 0 1 5076
box -55 -228 56 228
use M2_M1$$34864172_3v256x8m81  M2_M1$$34864172_3v256x8m81_0
timestamp 1763766357
transform 1 0 413 0 1 4570
box -119 -46 119 46
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_0
timestamp 1763766357
transform 1 0 339 0 1 1042
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_1
timestamp 1763766357
transform 1 0 645 0 1 2696
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_2
timestamp 1763766357
transform 1 0 1005 0 1 2696
box -43 -122 43 122
use M2_M1$$43377708_3v256x8m81  M2_M1$$43377708_3v256x8m81_0
timestamp 1763766357
transform 1 0 853 0 1 4005
box -44 -427 44 427
use M2_M1$$43377708_3v256x8m81  M2_M1$$43377708_3v256x8m81_1
timestamp 1763766357
transform 1 0 493 0 1 4005
box -44 -427 44 427
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_0
timestamp 1763766357
transform 1 0 339 0 1 5196
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_1
timestamp 1763766357
transform 1 0 484 0 1 5196
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_2
timestamp 1763766357
transform 1 0 848 0 1 5196
box -44 -275 44 275
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_0
timestamp 1763766357
transform 1 0 1188 0 1 2867
box -44 -123 44 123
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_1
timestamp 1763766357
transform 1 0 845 0 1 2534
box -44 -123 44 123
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_0
timestamp 1763766357
transform 1 0 339 0 1 5196
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_1
timestamp 1763766357
transform 1 0 484 0 1 5196
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_2
timestamp 1763766357
transform 1 0 848 0 1 5196
box -84 -185 84 275
use M3_M2$$47334444_3v256x8m81  M3_M2$$47334444_3v256x8m81_0
timestamp 1763766357
transform 1 0 853 0 1 4005
box -45 -427 45 427
use M3_M2$$47334444_3v256x8m81  M3_M2$$47334444_3v256x8m81_1
timestamp 1763766357
transform 1 0 493 0 1 4005
box -45 -427 45 427
use nmos_1p2$$47514668_3v256x8m81  nmos_1p2$$47514668_3v256x8m81_0
timestamp 1763766357
transform 1 0 907 0 1 4669
box -102 -44 130 467
use nmos_1p2$$47514668_3v256x8m81  nmos_1p2$$47514668_3v256x8m81_1
timestamp 1763766357
transform 1 0 547 0 1 4669
box -102 -44 130 467
use pmos_1p2$$46887980_3v256x8m81  pmos_1p2$$46887980_3v256x8m81_0
timestamp 1764700137
transform 1 0 907 0 1 2567
box -188 -86 216 1356
use pmos_1p2$$46887980_3v256x8m81  pmos_1p2$$46887980_3v256x8m81_1
timestamp 1764700137
transform 1 0 547 0 1 2567
box -188 -86 216 1356
<< end >>
