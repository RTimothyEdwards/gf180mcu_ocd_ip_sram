magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< nwell >>
rect -273 -154 273 154
<< nsubdiff >>
rect -170 23 170 54
rect -170 -23 -137 23
rect 137 -23 170 23
rect -170 -53 170 -23
<< nsubdiffcont >>
rect -137 -23 137 23
<< metal1 >>
rect -156 23 156 40
rect -156 -23 -137 23
rect 137 -23 156 23
rect -156 -39 156 -23
<< end >>
