magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< psubdiff >>
rect -1605 57 -1493 58
rect 1383 57 1605 58
rect -1605 23 1605 57
rect -1605 -23 -1351 23
rect 1351 -23 1605 23
rect -1605 -58 1605 -23
<< psubdiffcont >>
rect -1351 -23 1351 23
<< metal1 >>
rect -1599 23 1599 51
rect -1599 -23 -1351 23
rect 1351 -23 1599 23
rect -1599 -51 1599 -23
<< end >>
