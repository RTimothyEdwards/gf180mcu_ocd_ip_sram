magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< nwell >>
rect 1189 1215 1235 1833
<< polysilicon >>
rect 533 4306 589 5317
rect 893 4306 949 5321
<< metal1 >>
rect 227 5323 529 5964
rect 605 5337 686 5442
rect 605 5263 689 5337
rect 605 5179 901 5263
rect 245 3566 529 5026
rect 605 4149 686 5179
rect 965 4178 1045 5469
rect -74 3446 1276 3511
rect -74 3305 1276 3370
rect -74 3164 1276 3229
rect -74 3023 1276 3088
rect -74 2881 1276 2946
rect -74 2740 1276 2805
<< metal2 >>
rect 133 5364 526 5913
rect 736 5567 893 5913
rect 891 5552 893 5567
rect 133 5335 222 5364
rect 133 5110 221 5335
rect 294 1901 385 5178
rect 800 1879 890 3183
rect 1143 2230 1233 3374
rect 800 1786 1233 1879
<< metal3 >>
rect 0 5003 1276 5579
rect 0 3424 1184 4907
rect 4 3221 1233 3314
rect 9 2964 1270 3057
rect 800 2911 890 2964
use alatch_3v512x8m81  alatch_3v512x8m81_0
timestamp 1763765945
transform 1 0 49 0 1 443
box -63 409 1197 2033
use M1_NWELL10_3v512x8m81  M1_NWELL10_3v512x8m81_0
timestamp 1763765945
transform 1 0 233 0 1 4019
box -154 -530 154 1130
use M1_POLY2$$46559276_3v512x8m81  M1_POLY2$$46559276_3v512x8m81_0
timestamp 1763765945
transform 1 0 805 0 1 5221
box -123 -48 123 48
use M1_POLY2$$46559276_3v512x8m81  M1_POLY2$$46559276_3v512x8m81_1
timestamp 1763765945
transform 1 0 448 0 1 5221
box -123 -48 123 48
use M1_PSUB$$47335468_3v512x8m81  M1_PSUB$$47335468_3v512x8m81_0
timestamp 1763765945
transform 1 0 276 0 1 5537
box -55 -190 56 400
use M2_M1$$34864172_3v512x8m81  M2_M1$$34864172_3v512x8m81_0
timestamp 1763765945
transform 1 0 413 0 1 5221
box -119 -46 119 46
use M2_M1$$43375660_3v512x8m81  M2_M1$$43375660_3v512x8m81_0
timestamp 1763765945
transform 1 0 339 0 1 1042
box -43 -122 43 122
use M2_M1$$43375660_3v512x8m81  M2_M1$$43375660_3v512x8m81_1
timestamp 1763765945
transform 1 0 645 0 1 3696
box -43 -122 43 122
use M2_M1$$43375660_3v512x8m81  M2_M1$$43375660_3v512x8m81_2
timestamp 1763765945
transform 1 0 1005 0 1 3696
box -43 -122 43 122
use M2_M1$$43377708_3v512x8m81  M2_M1$$43377708_3v512x8m81_0
timestamp 1763765945
transform 1 0 853 0 1 4509
box -44 -427 44 427
use M2_M1$$43377708_3v512x8m81  M2_M1$$43377708_3v512x8m81_1
timestamp 1763765945
transform 1 0 493 0 1 4509
box -44 -427 44 427
use M2_M1$$43379756_3v512x8m81  M2_M1$$43379756_3v512x8m81_0
timestamp 1763765945
transform 1 0 339 0 1 5638
box -44 -275 44 275
use M2_M1$$43379756_3v512x8m81  M2_M1$$43379756_3v512x8m81_1
timestamp 1763765945
transform 1 0 484 0 1 5638
box -44 -275 44 275
use M2_M1$$43379756_3v512x8m81  M2_M1$$43379756_3v512x8m81_2
timestamp 1763765945
transform 1 0 848 0 1 5638
box -44 -275 44 275
use M2_M1_154_3v512x8m81  M2_M1_154_3v512x8m81_5
timestamp 1763765945
transform 1 0 339 0 1 1938
box -44 -123 44 122
use M3_M2$$43368492_3v512x8m81  M3_M2$$43368492_3v512x8m81_0
timestamp 1763765945
transform 1 0 1188 0 1 3237
box -44 -123 44 123
use M3_M2$$43368492_3v512x8m81  M3_M2$$43368492_3v512x8m81_1
timestamp 1763765945
transform 1 0 845 0 1 3034
box -44 -123 44 123
use M3_M2$$47333420_3v512x8m81  M3_M2$$47333420_3v512x8m81_0
timestamp 1763765945
transform 1 0 177 0 1 5294
box -84 -185 84 275
use M3_M2$$47333420_3v512x8m81  M3_M2$$47333420_3v512x8m81_1
timestamp 1763765945
transform 1 0 780 0 1 5306
box -84 -185 84 275
use M3_M2$$47334444_3v512x8m81  M3_M2$$47334444_3v512x8m81_0
timestamp 1763765945
transform 1 0 853 0 1 4469
box -45 -427 45 427
use M3_M2$$47334444_3v512x8m81  M3_M2$$47334444_3v512x8m81_1
timestamp 1763765945
transform 1 0 493 0 1 4469
box -45 -427 45 427
use nmos_1p2$$47336492_3v512x8m81  nmos_1p2$$47336492_3v512x8m81_0
timestamp 1763765945
transform 1 0 907 0 1 5349
box -102 -44 130 658
use nmos_1p2$$47336492_3v512x8m81  nmos_1p2$$47336492_3v512x8m81_1
timestamp 1763765945
transform 1 0 547 0 1 5349
box -102 -44 130 658
use pmos_1p2$$47337516_3v512x8m81  pmos_1p2$$47337516_3v512x8m81_0
timestamp 1763765945
transform 1 0 907 0 1 3567
box -188 -86 216 1610
use pmos_1p2$$47337516_3v512x8m81  pmos_1p2$$47337516_3v512x8m81_1
timestamp 1763765945
transform 1 0 547 0 1 3567
box -188 -86 216 1610
<< end >>
