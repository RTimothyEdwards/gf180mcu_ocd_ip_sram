magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal1 >>
rect -113 1146 113 1155
rect -113 -646 -105 1146
rect 105 -646 113 1146
rect -113 -655 113 -646
<< via1 >>
rect -105 -646 105 1146
<< metal2 >>
rect -113 1146 113 1155
rect -113 -646 -105 1146
rect 105 -646 113 1146
rect -113 -655 113 -646
<< end >>
