magic
tech gf180mcuD
magscale 1 10
timestamp 1763486358
<< nwell >>
rect -161 5039 54 8484
rect -121 1503 3715 2318
rect -121 642 3694 1503
<< metal1 >>
rect -16 6908 3476 6960
<< metal2 >>
rect 752 1055 814 1273
rect 1689 1055 1750 1267
rect 2591 1055 2652 1259
<< metal3 >>
rect -575 5420 4956 5618
use M1_NACTIVE4310591302028_512x8m81  M1_NACTIVE4310591302028_512x8m81_0
timestamp 1763476864
transform 1 0 426 0 1 5519
box -36 -95 36 95
use M1_NACTIVE4310591302028_512x8m81  M1_NACTIVE4310591302028_512x8m81_1
timestamp 1763476864
transform 1 0 1332 0 1 5519
box -36 -95 36 95
use M1_NACTIVE4310591302028_512x8m81  M1_NACTIVE4310591302028_512x8m81_2
timestamp 1763476864
transform 1 0 2236 0 1 5519
box -36 -95 36 95
use M1_NACTIVE4310591302028_512x8m81  M1_NACTIVE4310591302028_512x8m81_3
timestamp 1763476864
transform 1 0 3140 0 1 5519
box -36 -95 36 95
use M1_PACTIVE4310591302027_512x8m81  M1_PACTIVE4310591302027_512x8m81_0
timestamp 1763476864
transform 1 0 882 0 1 347
box -36 -62 36 62
use M1_PACTIVE4310591302027_512x8m81  M1_PACTIVE4310591302027_512x8m81_1
timestamp 1763476864
transform 1 0 1789 0 1 347
box -36 -62 36 62
use M1_PACTIVE4310591302027_512x8m81  M1_PACTIVE4310591302027_512x8m81_2
timestamp 1763476864
transform 1 0 3523 0 1 347
box -36 -62 36 62
use M1_PACTIVE4310591302027_512x8m81  M1_PACTIVE4310591302027_512x8m81_3
timestamp 1763476864
transform 1 0 2686 0 1 347
box -36 -62 36 62
use M1_PACTIVE4310591302027_512x8m81  M1_PACTIVE4310591302027_512x8m81_4
timestamp 1763476864
transform 1 0 -6 0 1 347
box -36 -62 36 62
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_0
timestamp 1763476864
transform 1 0 426 0 1 5519
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_1
timestamp 1763476864
transform 1 0 1332 0 1 5519
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_2
timestamp 1763476864
transform 1 0 2236 0 1 5519
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_3
timestamp 1763476864
transform 1 0 3140 0 1 5519
box -34 -99 34 99
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_2
timestamp 1763476864
transform 1 0 1719 0 1 1248
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_4
timestamp 1763476864
transform 1 0 2621 0 1 1248
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_5
timestamp 1763476864
transform 1 0 779 0 1 1248
box -35 -56 35 55
use M3_M2431059130201_512x8m81  M3_M2431059130201_512x8m81_1
timestamp 1763476864
transform 1 0 1719 0 1 1181
box -35 -63 35 63
use M3_M2431059130201_512x8m81  M3_M2431059130201_512x8m81_3
timestamp 1763476864
transform 1 0 2621 0 1 1181
box -35 -63 35 63
use M3_M2431059130201_512x8m81  M3_M2431059130201_512x8m81_5
timestamp 1763476864
transform 1 0 779 0 1 1231
box -35 -63 35 63
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_0
timestamp 1763476864
transform 1 0 426 0 1 5519
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_1
timestamp 1763476864
transform 1 0 1332 0 1 5519
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_2
timestamp 1763476864
transform 1 0 2236 0 1 5519
box -35 -99 35 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_3
timestamp 1763476864
transform 1 0 3140 0 1 5519
box -35 -99 35 99
use ypass_gate_512x8m81  ypass_gate_512x8m81_1
timestamp 1763485967
transform -1 0 3190 0 1 -3377
box -130 3470 633 11861
use ypass_gate_512x8m81  ypass_gate_512x8m81_2
timestamp 1763485967
transform -1 0 2288 0 1 -3377
box -130 3470 633 11861
use ypass_gate_512x8m81  ypass_gate_512x8m81_3
timestamp 1763485967
transform -1 0 1386 0 1 -3377
box -130 3470 633 11861
use ypass_gate_512x8m81  ypass_gate_512x8m81_4
timestamp 1763485967
transform 1 0 2180 0 1 -3377
box -130 3470 633 11861
use ypass_gate_512x8m81  ypass_gate_512x8m81_5
timestamp 1763485967
transform 1 0 1278 0 1 -3377
box -130 3470 633 11861
use ypass_gate_512x8m81  ypass_gate_512x8m81_6
timestamp 1763485967
transform 1 0 376 0 1 -3377
box -130 3470 633 11861
use ypass_gate_512x8m81  ypass_gate_512x8m81_7
timestamp 1763485967
transform -1 0 484 0 1 -3377
box -130 3470 633 11861
use ypass_gate_a_512x8m81  ypass_gate_a_512x8m81_0
timestamp 1763485967
transform 1 0 3090 0 1 -3377
box -130 3470 627 11860
<< end >>
