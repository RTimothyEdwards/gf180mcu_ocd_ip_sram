magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -70 410 70 417
rect -70 -410 -63 410
rect 63 -410 70 410
rect -70 -417 70 -410
<< via2 >>
rect -63 -410 63 410
<< metal3 >>
rect -70 410 70 417
rect -70 -410 -63 410
rect 63 -410 70 410
rect -70 -417 70 -410
<< end >>
