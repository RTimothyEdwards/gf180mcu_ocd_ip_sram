magic
tech gf180mcuD
magscale 1 10
timestamp 1765926640
<< nwell >>
rect -365 21493 15173 21547
rect 7182 21393 7401 21493
rect 14949 21393 15173 21493
rect -363 18111 15173 21393
rect 7571 18056 15173 18111
rect -363 14112 15178 14975
rect 3305 7222 3364 7239
rect 11073 7222 11116 7229
<< metal1 >>
rect 10403 12879 10675 12976
rect 10973 12879 11379 12976
rect -275 535 -44 587
rect 7037 533 7093 585
rect 7491 533 7547 585
rect 14808 533 14859 585
<< metal2 >>
rect -699 20267 -629 22826
rect -417 20264 -347 22826
rect 7116 20485 7186 22826
rect 7399 20491 7469 22826
rect 14931 20430 15001 22826
rect 15213 20448 15283 22826
<< metal3 >>
rect -771 99977 15976 100229
rect -771 99311 15976 99563
rect -771 98765 15976 99017
rect -771 98099 15976 98351
rect -771 97553 15976 97805
rect -771 96887 15976 97139
rect -771 96341 15976 96593
rect -771 95675 15976 95927
rect -771 95129 15976 95381
rect -771 94463 15976 94715
rect -771 93917 15976 94169
rect -771 93251 15976 93503
rect -771 92705 15976 92957
rect -771 92039 15976 92291
rect -771 91493 15976 91745
rect -771 90827 15976 91079
rect -771 90281 15976 90533
rect -771 89615 15976 89867
rect -771 89069 15976 89321
rect -771 88403 15976 88655
rect -771 87857 15976 88109
rect -771 87191 15976 87443
rect -771 86645 15976 86897
rect -771 85979 15976 86231
rect -771 85433 15976 85685
rect -771 84767 15976 85019
rect -771 84221 15976 84473
rect -771 83555 15976 83807
rect -771 83009 15976 83261
rect -771 82343 15976 82595
rect -771 81797 15976 82049
rect -771 81131 15976 81383
rect -771 80585 15976 80837
rect -771 79919 15976 80171
rect -771 79373 15976 79625
rect -771 78707 15976 78959
rect -771 78161 15976 78413
rect -771 77495 15976 77747
rect -771 76949 15976 77201
rect -771 76283 15976 76535
rect -771 75737 15976 75989
rect -771 75071 15976 75323
rect -771 74525 15976 74777
rect -771 73859 15976 74111
rect -771 73313 15976 73565
rect -771 72647 15976 72899
rect -771 72101 15976 72353
rect -771 71435 15976 71687
rect -771 70889 15976 71141
rect -771 70223 15976 70475
rect -771 69677 15976 69929
rect -771 69011 15976 69263
rect -771 68465 15976 68717
rect -771 67799 15976 68051
rect -771 67253 15976 67505
rect -771 66587 15976 66839
rect -771 66041 15976 66293
rect -771 65375 15976 65627
rect -771 64829 15976 65081
rect -771 64163 15976 64415
rect -771 63617 15976 63869
rect -771 62951 15976 63203
rect -771 62405 15976 62657
rect -771 61739 15976 61991
rect -771 61193 15976 61445
rect -771 60527 15976 60779
rect -771 59981 15976 60233
rect -771 59315 15976 59567
rect -771 58769 15976 59021
rect -771 58103 15976 58355
rect -771 57557 15976 57809
rect -771 56891 15976 57143
rect -771 56345 15976 56597
rect -771 55679 15976 55931
rect -771 55133 15976 55385
rect -771 54467 15976 54719
rect -771 53921 15976 54173
rect -771 53255 15976 53507
rect -771 52709 15976 52961
rect -771 52043 15976 52295
rect -771 51497 15976 51749
rect -771 50831 15976 51083
rect -771 50285 15976 50537
rect -771 49619 15976 49871
rect -771 49073 15976 49325
rect -771 48407 15976 48659
rect -771 47861 15976 48113
rect -771 47195 15976 47447
rect -771 46649 15976 46901
rect -771 45983 15976 46235
rect -771 45437 15976 45689
rect -771 44771 15976 45023
rect -771 44225 15976 44477
rect -771 43559 15976 43811
rect -771 43013 15976 43265
rect -771 42347 15976 42599
rect -771 41801 15976 42053
rect -771 41135 15976 41387
rect -771 40589 15976 40841
rect -771 39923 15976 40175
rect -771 39377 15976 39629
rect -771 38711 15976 38963
rect -771 38165 15976 38417
rect -771 37499 15976 37751
rect -771 36953 15976 37205
rect -771 36287 15976 36539
rect -771 35741 15976 35993
rect -771 35075 15976 35327
rect -771 34529 15976 34781
rect -771 33863 15976 34115
rect -771 33317 15976 33569
rect -771 32651 15976 32903
rect -771 32105 15976 32357
rect -771 31439 15976 31691
rect -771 30893 15976 31145
rect -771 30227 15976 30479
rect -771 29681 15976 29933
rect -771 29015 15976 29267
rect -771 28469 15976 28721
rect -771 27803 15976 28055
rect -771 27257 15976 27509
rect -771 26591 15976 26843
rect -771 26045 15976 26297
rect -771 25379 15976 25631
rect -771 24833 15976 25085
rect -771 24167 15976 24419
rect -771 23621 15976 23873
rect -771 22955 15976 23207
rect -771 22409 15976 22661
rect -821 21665 15523 22001
rect -821 20111 15523 21377
rect -461 16504 14939 16654
rect -461 16265 14939 16416
rect -461 16021 14939 16171
rect -461 15780 14939 15931
rect -461 15553 14939 15703
rect -461 15307 14939 15458
rect -461 15063 14939 15213
rect -461 14817 14939 14968
rect -461 14363 14939 14672
rect -461 13648 14939 13967
rect -461 11041 14939 12947
rect -461 10047 14539 10840
rect -461 8983 14939 10047
rect -481 8356 14939 8858
rect -481 7425 14939 7992
rect -461 6121 14939 7043
rect 659 6018 13680 6021
rect -124 5960 13680 6018
rect -461 4706 14939 5660
rect -461 4125 14939 4489
rect -461 3720 14939 4061
rect -461 3355 14939 3657
rect -461 2940 14939 3259
rect -487 2238 15003 2557
rect -487 1792 15003 2037
rect -487 1644 15003 1705
rect -487 1481 15003 1542
rect -487 1149 15003 1394
rect -487 641 15003 960
use Cell_array8x8_3v1024x8m81  Cell_array8x8_3v1024x8m81_0
timestamp 1765925964
transform 1 0 -996 0 1 22638
box 262 103 16314 77801
use M3_M24310591302022_3v1024x8m81  M3_M24310591302022_3v1024x8m81_0
timestamp 1764525316
transform 1 0 14966 0 1 20765
box -35 -534 35 534
use M3_M24310591302022_3v1024x8m81  M3_M24310591302022_3v1024x8m81_1
timestamp 1764525316
transform 1 0 -379 0 1 20825
box -35 -534 35 534
use M3_M24310591302022_3v1024x8m81  M3_M24310591302022_3v1024x8m81_2
timestamp 1764525316
transform 1 0 7430 0 1 20825
box -35 -534 35 534
use M3_M24310591302023_3v1024x8m81  M3_M24310591302023_3v1024x8m81_0
timestamp 1764525316
transform 1 0 7152 0 1 21835
box -35 -165 35 165
use M3_M24310591302023_3v1024x8m81  M3_M24310591302023_3v1024x8m81_1
timestamp 1764525316
transform 1 0 -659 0 1 21835
box -35 -165 35 165
use M3_M24310591302023_3v1024x8m81  M3_M24310591302023_3v1024x8m81_2
timestamp 1764525316
transform 1 0 15250 0 1 21835
box -35 -165 35 165
use saout_m2_3v1024x8m81  saout_m2_3v1024x8m81_3
timestamp 1765925964
transform 1 0 -591 0 1 1002
box -188 -475 5343 21797
use saout_m2_3v1024x8m81  saout_m2_3v1024x8m81_4
timestamp 1765925964
transform 1 0 7175 0 1 1002
box -188 -475 5343 21797
use saout_R_m2_3v1024x8m81  saout_R_m2_3v1024x8m81_0
timestamp 1765925964
transform -1 0 15175 0 1 1007
box -188 -482 5343 21793
use saout_R_m2_3v1024x8m81  saout_R_m2_3v1024x8m81_1
timestamp 1765925964
transform -1 0 7409 0 1 1007
box -188 -482 5343 21793
<< labels >>
flabel metal3 s -219 21842 -219 21842 0 FreeSans 313 0 0 0 VSS
port 76 nsew
flabel metal3 s -219 17082 -219 17082 0 FreeSans 313 0 0 0 VSS
port 76 nsew
rlabel metal2 s -159 21313 -159 21313 4 b[31]
port 87 nsew
rlabel metal2 s 707 21313 707 21313 4 b[29]
port 96 nsew
rlabel metal2 s 273 21313 273 21313 4 bb[30]
port 136 nsew
rlabel metal1 s 11515 12152 11515 12152 4 pcb[0]
port 149 nsew
rlabel metal1 s 9965 12152 9965 12152 4 pcb[1]
port 150 nsew
rlabel metal1 s 2579 12152 2579 12152 4 pcb[3]
port 151 nsew
rlabel metal1 s 3939 12152 3939 12152 4 pcb[2]
port 152 nsew
rlabel metal3 s -500 23132 -500 23132 4 WL[0]
port 72 nsew
rlabel metal3 s -500 23714 -500 23714 4 WL[1]
port 12 nsew
rlabel metal3 s -500 24344 -500 24344 4 WL[2]
port 11 nsew
rlabel metal3 s -500 24926 -500 24926 4 WL[3]
port 1 nsew
rlabel metal3 s -500 25556 -500 25556 4 WL[4]
port 52 nsew
rlabel metal3 s -500 26138 -500 26138 4 WL[5]
port 49 nsew
rlabel metal3 s -500 26768 -500 26768 4 WL[6]
port 46 nsew
rlabel metal3 s -500 27980 -500 27980 4 WL[8]
port 41 nsew
rlabel metal3 s -500 27350 -500 27350 4 WL[7]
port 44 nsew
rlabel metal3 s -500 28562 -500 28562 4 WL[9]
port 36 nsew
rlabel metal3 s -500 29192 -500 29192 4 WL[10]
port 35 nsew
rlabel metal3 s -500 29774 -500 29774 4 WL[11]
port 30 nsew
rlabel metal3 s -500 30404 -500 30404 4 WL[12]
port 29 nsew
rlabel metal3 s -500 30986 -500 30986 4 WL[13]
port 68 nsew
rlabel metal3 s -500 31616 -500 31616 4 WL[14]
port 65 nsew
rlabel metal3 s -500 32198 -500 32198 4 WL[15]
port 64 nsew
rlabel metal3 s -500 32828 -500 32828 4 WL[16]
port 61 nsew
rlabel metal3 s -500 33410 -500 33410 4 WL[17]
port 58 nsew
rlabel metal3 s -500 34040 -500 34040 4 WL[18]
port 55 nsew
rlabel metal3 s -500 34622 -500 34622 4 WL[19]
port 24 nsew
rlabel metal3 s -500 35252 -500 35252 4 WL[20]
port 23 nsew
rlabel metal3 s -500 36464 -500 36464 4 WL[22]
port 19 nsew
rlabel metal3 s -500 35834 -500 35834 4 WL[21]
port 20 nsew
rlabel metal3 s -500 37046 -500 37046 4 WL[23]
port 18 nsew
rlabel metal3 s -500 37676 -500 37676 4 WL[24]
port 17 nsew
rlabel metal3 s -500 38258 -500 38258 4 WL[25]
port 75 nsew
rlabel metal3 s -500 38888 -500 38888 4 WL[26]
port 71 nsew
rlabel metal3 s -500 39470 -500 39470 4 WL[27]
port 70 nsew
rlabel metal3 s -500 40100 -500 40100 4 WL[28]
port 69 nsew
rlabel metal3 s -500 40682 -500 40682 4 WL[29]
port 16 nsew
rlabel metal3 s -500 41312 -500 41312 4 WL[30]
port 15 nsew
rlabel metal3 s -500 41894 -500 41894 4 WL[31]
port 14 nsew
rlabel metal3 s -500 42522 -500 42522 4 WL[32]
port 13 nsew
rlabel metal3 s -500 43104 -500 43104 4 WL[33]
port 45 nsew
rlabel metal3 s -500 43734 -500 43734 4 WL[34]
port 40 nsew
rlabel metal3 s -500 44316 -500 44316 4 WL[35]
port 39 nsew
rlabel metal3 s -500 44946 -500 44946 4 WL[36]
port 48 nsew
rlabel metal3 s -500 45528 -500 45528 4 WL[37]
port 43 nsew
rlabel metal3 s -500 46158 -500 46158 4 WL[38]
port 47 nsew
rlabel metal3 s -500 46740 -500 46740 4 WL[39]
port 42 nsew
rlabel metal3 s -500 47370 -500 47370 4 WL[40]
port 34 nsew
rlabel metal3 s -500 47952 -500 47952 4 WL[41]
port 33 nsew
rlabel metal3 s -500 48582 -500 48582 4 WL[42]
port 37 nsew
rlabel metal3 s -500 49164 -500 49164 4 WL[43]
port 38 nsew
rlabel metal3 s -500 49794 -500 49794 4 WL[44]
port 54 nsew
rlabel metal3 s -500 50376 -500 50376 4 WL[45]
port 51 nsew
rlabel metal3 s -500 51006 -500 51006 4 WL[46]
port 53 nsew
rlabel metal3 s -500 51588 -500 51588 4 WL[47]
port 50 nsew
rlabel metal3 s -500 52223 -500 52223 4 WL[48]
port 28 nsew
rlabel metal3 s -500 52805 -500 52805 4 WL[49]
port 27 nsew
rlabel metal3 s -500 53435 -500 53435 4 WL[50]
port 31 nsew
rlabel metal3 s -500 54017 -500 54017 4 WL[51]
port 32 nsew
rlabel metal3 s -500 54647 -500 54647 4 WL[52]
port 60 nsew
rlabel metal3 s -500 55229 -500 55229 4 WL[53]
port 57 nsew
rlabel metal3 s -500 55859 -500 55859 4 WL[54]
port 59 nsew
rlabel metal3 s -500 56441 -500 56441 4 WL[55]
port 56 nsew
rlabel metal3 s -500 57071 -500 57071 4 WL[56]
port 22 nsew
rlabel metal3 s -500 57653 -500 57653 4 WL[57]
port 21 nsew
rlabel metal3 s -500 58283 -500 58283 4 WL[58]
port 25 nsew
rlabel metal3 s -500 58865 -500 58865 4 WL[59]
port 26 nsew
rlabel metal3 s -500 59495 -500 59495 4 WL[60]
port 67 nsew
rlabel metal3 s -500 60077 -500 60077 4 WL[61]
port 63 nsew
rlabel metal3 s -500 60707 -500 60707 4 WL[62]
port 66 nsew
rlabel metal2 s 10738 21313 10738 21313 4 bb[8]
port 114 nsew
rlabel metal2 s 9871 21313 9871 21313 4 bb[10]
port 116 nsew
rlabel metal2 s 9729 21313 9729 21313 4 bb[11]
port 117 nsew
rlabel metal2 s 9296 21313 9296 21313 4 b[12]
port 142 nsew
rlabel metal2 s 10304 21313 10304 21313 4 b[9]
port 143 nsew
flabel metal3 s -219 20551 -219 20551 0 FreeSans 313 0 0 0 VDD
port 10 nsew
rlabel metal3 s 567 15835 567 15835 4 ypass[4]
port 5 nsew
rlabel metal3 s 567 16077 567 16077 4 ypass[5]
port 6 nsew
rlabel metal3 s 567 16318 567 16318 4 ypass[6]
port 73 nsew
rlabel metal3 s 567 16554 567 16554 4 ypass[7]
port 7 nsew
rlabel metal3 s 567 15633 567 15633 4 ypass[3]
port 4 nsew
rlabel metal3 s 567 15391 567 15391 4 ypass[2]
port 74 nsew
rlabel metal3 s 567 15149 567 15149 4 ypass[1]
port 3 nsew
rlabel metal3 s 567 14903 567 14903 4 ypass[0]
port 2 nsew
flabel metal3 s -219 14516 -219 14516 0 FreeSans 313 0 0 0 VDD
port 10 nsew
flabel metal3 s -219 13853 -219 13853 0 FreeSans 313 0 0 0 VSS
port 76 nsew
flabel metal3 s -219 9967 -219 9967 0 FreeSans 313 0 0 0 VSS
port 76 nsew
flabel metal3 s -219 11750 -219 11750 0 FreeSans 313 0 0 0 VDD
port 10 nsew
flabel metal3 s -219 7820 -219 7820 0 FreeSans 313 0 0 0 VDD
port 10 nsew
flabel metal3 s -219 6659 -219 6659 0 FreeSans 313 0 0 0 VSS
port 76 nsew
flabel metal3 s -219 5214 -219 5214 0 FreeSans 313 0 0 0 VDD
port 10 nsew
flabel metal3 s -219 4313 -219 4313 0 FreeSans 313 0 0 0 VSS
port 76 nsew
rlabel metal3 s 616 3790 616 3790 4 men
port 8 nsew
flabel metal3 s -219 3530 -219 3530 0 FreeSans 313 0 0 0 VSS
port 76 nsew
flabel metal3 s -219 3105 -219 3105 0 FreeSans 313 0 0 0 VDD
port 10 nsew
flabel metal3 s -219 2393 -219 2393 0 FreeSans 313 0 0 0 VDD
port 10 nsew
flabel metal3 s -219 774 -219 774 0 FreeSans 313 0 0 0 VDD
port 10 nsew
flabel metal1 s -247 562 -247 562 0 FreeSans 420 0 0 0 WEN[3]
port 153 nsew
flabel metal1 s 7057 558 7057 558 0 FreeSans 420 0 0 0 WEN[2]
port 154 nsew
flabel metal1 s 7514 558 7514 558 0 FreeSans 420 0 0 0 WEN[1]
port 155 nsew
flabel metal1 s 14832 558 14832 558 0 FreeSans 420 0 0 0 WEN[0]
port 156 nsew
flabel metal3 s -109 5987 -109 5987 0 FreeSans 313 0 0 0 GWE
port 9 nsew
rlabel metal3 s -500 100073 -500 100073 4 WL[127]
port 62 nsew
rlabel metal2 s -240 2832 -240 2832 4 din[0]
port 91 nsew
rlabel metal2 s 402 2888 402 2888 4 q[0]
port 92 nsew
rlabel metal2 s 6447 2928 6447 2928 4 q[1]
port 93 nsew
rlabel metal2 s 7049 2951 7049 2951 4 din[1]
port 88 nsew
rlabel metal2 s 7536 2832 7536 2832 4 din[2]
port 90 nsew
rlabel metal2 s 8148 2888 8148 2888 4 q[2]
port 94 nsew
rlabel metal2 s 14199 2925 14199 2925 4 q[3]
port 95 nsew
rlabel metal2 s 14818 2949 14818 2949 4 din[3]
port 89 nsew
rlabel metal2 s 162 21313 162 21313 4 bb[31]
port 137 nsew
rlabel metal2 s 616 21303 616 21303 4 b[30]
port 138 nsew
rlabel metal2 s 1059 21313 1059 21313 4 bb[29]
port 135 nsew
rlabel metal2 s 1191 21313 1191 21313 4 bb[28]
port 134 nsew
rlabel metal2 s 1522 21313 1522 21313 4 b[28]
port 86 nsew
rlabel metal2 s 1634 21303 1634 21303 4 b[27]
port 139 nsew
rlabel metal2 s 1966 21323 1966 21323 4 bb[27]
port 133 nsew
rlabel metal2 s 2098 21323 2098 21323 4 bb[26]
port 132 nsew
rlabel metal2 s 6985 21313 6985 21313 4 b[16]
port 82 nsew
rlabel metal2 s 6652 21313 6652 21313 4 bb[16]
port 122 nsew
rlabel metal2 s 6531 21313 6531 21313 4 bb[17]
port 123 nsew
rlabel metal2 s 6189 21303 6189 21303 4 b[17]
port 100 nsew
rlabel metal2 s 6088 21313 6088 21313 4 b[18]
port 148 nsew
rlabel metal2 s 5756 21313 5756 21313 4 bb[18]
port 124 nsew
rlabel metal2 s 5624 21313 5624 21313 4 bb[19]
port 125 nsew
rlabel metal2 s 5302 21313 5302 21313 4 b[19]
port 83 nsew
rlabel metal2 s 5190 21313 5190 21313 4 b[20]
port 99 nsew
rlabel metal2 s 4848 21323 4848 21323 4 bb[20]
port 126 nsew
rlabel metal2 s 4727 21323 4727 21323 4 bb[21]
port 127 nsew
rlabel metal2 s 4395 21313 4395 21313 4 b[21]
port 144 nsew
rlabel metal2 s 4284 21313 4284 21313 4 b[22]
port 84 nsew
rlabel metal2 s 3952 21323 3952 21323 4 bb[22]
port 128 nsew
rlabel metal2 s 3830 21323 3830 21323 4 bb[23]
port 129 nsew
rlabel metal2 s 3468 21313 3468 21313 4 b[23]
port 98 nsew
rlabel metal2 s 3356 21323 3356 21323 4 b[24]
port 140 nsew
rlabel metal2 s 2994 21323 2994 21323 4 bb[24]
port 130 nsew
rlabel metal2 s 2873 21323 2873 21323 4 bb[25]
port 131 nsew
rlabel metal2 s 2541 21313 2541 21313 4 b[25]
port 85 nsew
rlabel metal2 s 2430 21313 2430 21313 4 b[26]
port 97 nsew
rlabel metal2 s 7593 21323 7593 21323 4 b[15]
port 141 nsew
rlabel metal2 s 7925 21323 7925 21323 4 bb[15]
port 121 nsew
rlabel metal2 s 8057 21313 8057 21313 4 bb[14]
port 120 nsew
rlabel metal2 s 8399 21313 8399 21313 4 b[14]
port 101 nsew
rlabel metal2 s 8510 21313 8510 21313 4 b[13]
port 81 nsew
rlabel metal2 s 8843 21303 8843 21303 4 bb[13]
port 119 nsew
rlabel metal2 s 8964 21313 8964 21313 4 bb[12]
port 118 nsew
rlabel metal2 s 9417 21323 9417 21323 4 b[11]
port 102 nsew
rlabel metal2 s 10193 21323 10193 21323 4 b[10]
port 80 nsew
rlabel metal2 s 10637 21313 10637 21313 4 bb[9]
port 115 nsew
rlabel metal2 s 11120 21323 11120 21323 4 b[8]
port 103 nsew
rlabel metal2 s 14758 21323 14758 21323 4 b[0]
port 145 nsew
rlabel metal2 s 14426 21323 14426 21323 4 bb[0]
port 106 nsew
rlabel metal2 s 14294 21323 14294 21323 4 bb[1]
port 107 nsew
rlabel metal2 s 13972 21323 13972 21323 4 b[1]
port 77 nsew
rlabel metal2 s 13851 21333 13851 21333 4 b[2]
port 105 nsew
rlabel metal2 s 13508 21333 13508 21333 4 bb[2]
port 108 nsew
rlabel metal2 s 13407 21323 13407 21323 4 bb[3]
port 109 nsew
rlabel metal2 s 13065 21333 13065 21333 4 b[3]
port 146 nsew
rlabel metal2 s 12954 21333 12954 21333 4 b[4]
port 78 nsew
rlabel metal2 s 12612 21323 12612 21323 4 bb[4]
port 110 nsew
rlabel metal2 s 12490 21333 12490 21333 4 bb[5]
port 111 nsew
rlabel metal2 s 12169 21323 12169 21323 4 b[5]
port 104 nsew
rlabel metal2 s 12047 21323 12047 21323 4 b[6]
port 147 nsew
rlabel metal2 s 11715 21333 11715 21333 4 bb[6]
port 112 nsew
rlabel metal2 s 11613 21333 11613 21333 4 bb[7]
port 113 nsew
rlabel metal2 s 11231 21313 11231 21313 4 b[7]
port 79 nsew
<< end >>
