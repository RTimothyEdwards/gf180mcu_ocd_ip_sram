magic
tech gf180mcuD
magscale 1 10
timestamp 1765833244
<< metal2 >>
rect -102 63 -33 1507
rect 111 186 181 1507
rect 335 352 405 1507
rect 547 458 617 1507
rect 547 388 659 458
rect 335 282 427 352
rect 111 116 303 186
rect -102 -6 -30 63
rect -86 -44 -30 -6
rect 247 -44 303 116
rect 371 -44 427 282
rect 589 192 659 388
rect 771 349 841 1507
rect 983 457 1053 1507
rect 983 387 1092 457
rect 771 279 872 349
rect 589 122 760 192
rect 704 -44 760 122
rect 816 -44 872 279
rect 1022 197 1092 387
rect 1207 341 1277 1507
rect 1419 460 1489 1507
rect 1419 390 1525 460
rect 1207 271 1329 341
rect 1022 127 1205 197
rect 1148 -44 1205 127
rect 1273 -44 1329 271
rect 1455 219 1525 390
rect 1643 362 1713 1507
rect 1643 292 1774 362
rect 1455 149 1662 219
rect 1606 -44 1662 149
rect 1718 -44 1774 292
rect 1855 213 1925 1507
rect 2078 354 2148 1507
rect 2078 284 2231 354
rect 1855 143 2107 213
rect 2051 -44 2107 143
rect 2175 -44 2231 284
rect 2291 197 2361 1507
rect 2515 345 2585 1507
rect 2727 485 2797 1507
rect 2727 415 2825 485
rect 2515 275 2676 345
rect 2291 127 2564 197
rect 2508 -44 2564 127
rect 2620 -44 2676 275
rect 2755 212 2825 415
rect 2951 341 3021 1507
rect 3163 482 3233 1507
rect 3163 412 3258 482
rect 2951 271 3121 341
rect 2755 142 3009 212
rect 2953 -44 3009 142
rect 3065 -44 3121 271
rect 3188 192 3258 412
rect 3188 122 3491 192
rect 3435 -44 3491 122
<< properties >>
string path 13.205 10.765 13.205 2.845 14.705 2.845 14.705 -0.315 
<< end >>
