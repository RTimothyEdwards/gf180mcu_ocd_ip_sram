magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal2 >>
rect -44 93 44 112
rect -44 -93 -28 93
rect 28 -93 44 93
rect -44 -111 44 -93
<< via2 >>
rect -28 -93 28 93
<< metal3 >>
rect -45 93 45 112
rect -45 -93 -28 93
rect 28 -93 45 93
rect -45 -112 45 -93
<< end >>
