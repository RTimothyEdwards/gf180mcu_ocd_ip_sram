magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nmos >>
rect -532 0 -476 687
rect -372 0 -316 687
rect -211 0 -155 687
rect -51 0 5 687
rect 110 0 166 687
rect 270 0 326 687
rect 431 0 487 687
rect 591 0 647 687
rect 752 0 808 687
rect 912 0 968 687
rect 1073 0 1129 687
rect 1233 0 1289 687
rect 1394 0 1450 687
rect 1554 0 1610 687
rect 1715 0 1771 687
rect 1876 0 1932 687
rect 2036 0 2092 687
rect 2197 0 2253 687
rect 2357 0 2413 687
rect 2518 0 2574 687
<< ndiff >>
rect -620 674 -532 687
rect -620 13 -607 674
rect -561 13 -532 674
rect -620 0 -532 13
rect -476 674 -372 687
rect -476 13 -447 674
rect -401 13 -372 674
rect -476 0 -372 13
rect -316 674 -211 687
rect -316 13 -286 674
rect -240 13 -211 674
rect -316 0 -211 13
rect -155 674 -51 687
rect -155 13 -126 674
rect -80 13 -51 674
rect -155 0 -51 13
rect 5 674 110 687
rect 5 13 34 674
rect 80 13 110 674
rect 5 0 110 13
rect 166 674 270 687
rect 166 13 195 674
rect 241 13 270 674
rect 166 0 270 13
rect 326 674 431 687
rect 326 13 355 674
rect 401 13 431 674
rect 326 0 431 13
rect 487 674 591 687
rect 487 13 516 674
rect 562 13 591 674
rect 487 0 591 13
rect 647 674 752 687
rect 647 13 676 674
rect 722 13 752 674
rect 647 0 752 13
rect 808 674 912 687
rect 808 13 837 674
rect 883 13 912 674
rect 808 0 912 13
rect 968 674 1073 687
rect 968 13 997 674
rect 1043 13 1073 674
rect 968 0 1073 13
rect 1129 674 1233 687
rect 1129 13 1158 674
rect 1204 13 1233 674
rect 1129 0 1233 13
rect 1289 674 1394 687
rect 1289 13 1318 674
rect 1364 13 1394 674
rect 1289 0 1394 13
rect 1450 674 1554 687
rect 1450 13 1479 674
rect 1525 13 1554 674
rect 1450 0 1554 13
rect 1610 674 1715 687
rect 1610 13 1639 674
rect 1685 13 1715 674
rect 1610 0 1715 13
rect 1771 674 1876 687
rect 1771 13 1800 674
rect 1846 13 1876 674
rect 1771 0 1876 13
rect 1932 674 2036 687
rect 1932 13 1961 674
rect 2007 13 2036 674
rect 1932 0 2036 13
rect 2092 674 2197 687
rect 2092 13 2121 674
rect 2167 13 2197 674
rect 2092 0 2197 13
rect 2253 674 2357 687
rect 2253 13 2282 674
rect 2328 13 2357 674
rect 2253 0 2357 13
rect 2413 674 2518 687
rect 2413 13 2442 674
rect 2488 13 2518 674
rect 2413 0 2518 13
rect 2574 674 2662 687
rect 2574 13 2603 674
rect 2649 13 2662 674
rect 2574 0 2662 13
<< ndiffc >>
rect -607 13 -561 674
rect -447 13 -401 674
rect -286 13 -240 674
rect -126 13 -80 674
rect 34 13 80 674
rect 195 13 241 674
rect 355 13 401 674
rect 516 13 562 674
rect 676 13 722 674
rect 837 13 883 674
rect 997 13 1043 674
rect 1158 13 1204 674
rect 1318 13 1364 674
rect 1479 13 1525 674
rect 1639 13 1685 674
rect 1800 13 1846 674
rect 1961 13 2007 674
rect 2121 13 2167 674
rect 2282 13 2328 674
rect 2442 13 2488 674
rect 2603 13 2649 674
<< polysilicon >>
rect -532 687 -476 731
rect -372 687 -316 731
rect -211 687 -155 731
rect -51 687 5 731
rect 110 687 166 731
rect 270 687 326 731
rect 431 687 487 731
rect 591 687 647 731
rect 752 687 808 731
rect 912 687 968 731
rect 1073 687 1129 731
rect 1233 687 1289 731
rect 1394 687 1450 731
rect 1554 687 1610 731
rect 1715 687 1771 731
rect 1876 687 1932 731
rect 2036 687 2092 731
rect 2197 687 2253 731
rect 2357 687 2413 731
rect 2518 687 2574 731
rect -532 -44 -476 0
rect -372 -44 -316 0
rect -211 -44 -155 0
rect -51 -44 5 0
rect 110 -44 166 0
rect 270 -44 326 0
rect 431 -44 487 0
rect 591 -44 647 0
rect 752 -44 808 0
rect 912 -44 968 0
rect 1073 -44 1129 0
rect 1233 -44 1289 0
rect 1394 -44 1450 0
rect 1554 -44 1610 0
rect 1715 -44 1771 0
rect 1876 -44 1932 0
rect 2036 -44 2092 0
rect 2197 -44 2253 0
rect 2357 -44 2413 0
rect 2518 -44 2574 0
<< metal1 >>
rect -607 674 -561 687
rect -607 0 -561 13
rect -447 674 -401 687
rect -447 0 -401 13
rect -286 674 -240 687
rect -286 0 -240 13
rect -126 674 -80 687
rect -126 0 -80 13
rect 34 674 80 687
rect 34 0 80 13
rect 195 674 241 687
rect 195 0 241 13
rect 355 674 401 687
rect 355 0 401 13
rect 516 674 562 687
rect 516 0 562 13
rect 676 674 722 687
rect 676 0 722 13
rect 837 674 883 687
rect 837 0 883 13
rect 997 674 1043 687
rect 997 0 1043 13
rect 1158 674 1204 687
rect 1158 0 1204 13
rect 1318 674 1364 687
rect 1318 0 1364 13
rect 1479 674 1525 687
rect 1479 0 1525 13
rect 1639 674 1685 687
rect 1639 0 1685 13
rect 1800 674 1846 687
rect 1800 0 1846 13
rect 1961 674 2007 687
rect 1961 0 2007 13
rect 2121 674 2167 687
rect 2121 0 2167 13
rect 2282 674 2328 687
rect 2282 0 2328 13
rect 2442 674 2488 687
rect 2442 0 2488 13
rect 2603 674 2649 687
rect 2603 0 2649 13
<< labels >>
flabel ndiffc 1021 343 1021 343 0 FreeSans 93 0 0 0 S
flabel ndiffc 872 343 872 343 0 FreeSans 93 0 0 0 D
flabel ndiffc 712 343 712 343 0 FreeSans 93 0 0 0 S
flabel ndiffc 551 343 551 343 0 FreeSans 93 0 0 0 D
flabel ndiffc 390 343 390 343 0 FreeSans 93 0 0 0 S
flabel ndiffc 230 343 230 343 0 FreeSans 93 0 0 0 D
flabel ndiffc 69 343 69 343 0 FreeSans 93 0 0 0 S
flabel ndiffc -91 343 -91 343 0 FreeSans 93 0 0 0 D
flabel ndiffc -252 343 -252 343 0 FreeSans 93 0 0 0 S
flabel ndiffc -412 343 -412 343 0 FreeSans 93 0 0 0 D
flabel ndiffc -572 343 -572 343 0 FreeSans 93 0 0 0 S
flabel ndiffc 1169 343 1169 343 0 FreeSans 93 0 0 0 D
flabel ndiffc 1330 343 1330 343 0 FreeSans 93 0 0 0 S
flabel ndiffc 1490 343 1490 343 0 FreeSans 93 0 0 0 D
flabel ndiffc 1651 343 1651 343 0 FreeSans 93 0 0 0 S
flabel ndiffc 1972 343 1972 343 0 FreeSans 93 0 0 0 S
flabel ndiffc 2132 343 2132 343 0 FreeSans 93 0 0 0 D
flabel ndiffc 2293 343 2293 343 0 FreeSans 93 0 0 0 S
flabel ndiffc 2614 343 2614 343 0 FreeSans 93 0 0 0 S
flabel ndiffc 2452 343 2452 343 0 FreeSans 93 0 0 0 D
flabel ndiffc 1810 343 1810 343 0 FreeSans 93 0 0 0 D
<< end >>
