magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal2 >>
rect -330 453 330 460
rect -330 -453 -323 453
rect 323 -453 330 453
rect -330 -460 330 -453
<< via2 >>
rect -323 -453 323 453
<< metal3 >>
rect -330 453 330 460
rect -330 -453 -323 453
rect 323 -453 330 453
rect -330 -460 330 -453
<< end >>
