magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< error_p >>
rect -79 -4 -33 64
rect 89 -3 135 65
<< nmos >>
rect 0 0 56 61
<< ndiff >>
rect -92 61 -20 66
rect 76 61 148 67
rect -92 53 0 61
rect -92 7 -79 53
rect -33 7 0 53
rect -92 0 0 7
rect 56 54 148 61
rect 56 8 89 54
rect 135 8 148 54
rect 56 0 148 8
rect -92 -6 -20 0
rect 76 -5 148 0
<< ndiffc >>
rect -79 7 -33 53
rect 89 8 135 54
<< polysilicon >>
rect 0 61 56 105
rect 0 -44 56 0
<< metal1 >>
rect -79 53 -33 64
rect -79 -4 -33 7
rect 89 54 135 65
rect 89 -3 135 8
<< labels >>
flabel ndiffc -44 30 -44 30 0 FreeSans 93 0 0 0 S
flabel ndiffc 100 30 100 30 0 FreeSans 93 0 0 0 D
<< end >>
