magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< psubdiff >>
rect -128 81 128 95
rect -128 -81 -114 81
rect 114 -81 128 81
rect -128 -95 128 -81
<< psubdiffcont >>
rect -114 -81 114 81
<< metal1 >>
rect -122 81 122 89
rect -122 -81 -114 81
rect 114 -81 122 81
rect -122 -89 122 -81
<< end >>
