magic
tech gf180mcuD
magscale 1 10
timestamp 1764700137
<< nmos >>
rect 0 0 56 635
<< ndiff >>
rect -88 622 0 635
rect -88 13 -75 622
rect -29 13 0 622
rect -88 0 0 13
rect 56 622 144 635
rect 56 13 85 622
rect 131 13 144 622
rect 56 0 144 13
<< ndiffc >>
rect -75 13 -29 622
rect 85 13 131 622
<< polysilicon >>
rect 0 635 56 679
rect 0 -44 56 0
<< metal1 >>
rect -75 622 -29 635
rect -75 0 -29 13
rect 85 622 131 635
rect 85 0 131 13
<< labels >>
flabel ndiffc -40 317 -40 317 0 FreeSans 93 0 0 0 S
flabel ndiffc 96 317 96 317 0 FreeSans 93 0 0 0 D
<< end >>
