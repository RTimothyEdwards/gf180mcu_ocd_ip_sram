magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< error_p >>
rect -103 0 -57 112
rect 57 0 103 112
rect 217 0 263 112
<< nmos >>
rect -28 0 28 112
rect 132 0 188 112
<< ndiff >>
rect -116 99 -28 112
rect -116 13 -103 99
rect -57 13 -28 99
rect -116 0 -28 13
rect 28 99 132 112
rect 28 13 57 99
rect 103 13 132 99
rect 28 0 132 13
rect 188 99 276 112
rect 188 13 217 99
rect 263 13 276 99
rect 188 0 276 13
<< ndiffc >>
rect -103 13 -57 99
rect 57 13 103 99
rect 217 13 263 99
<< polysilicon >>
rect -28 112 28 156
rect 132 112 188 156
rect -28 -44 28 0
rect 132 -44 188 0
<< metal1 >>
rect -103 99 -57 112
rect -103 0 -57 13
rect 57 99 103 112
rect 57 0 103 13
rect 217 99 263 112
rect 217 0 263 13
<< labels >>
flabel ndiffc 80 56 80 56 0 FreeSans 93 0 0 0 D
flabel ndiffc -68 56 -68 56 0 FreeSans 93 0 0 0 S
flabel ndiffc 228 56 228 56 0 FreeSans 93 0 0 0 S
<< end >>
