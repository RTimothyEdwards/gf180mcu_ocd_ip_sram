magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< psubdiff >>
rect -1328 73 1328 114
rect -1328 -73 -1288 73
rect 1288 -73 1328 73
rect -1328 -114 1328 -73
<< psubdiffcont >>
rect -1288 -73 1288 73
<< metal1 >>
rect -1323 73 1323 108
rect -1323 -73 -1288 73
rect 1288 -73 1323 73
rect -1323 -108 1323 -73
<< end >>
