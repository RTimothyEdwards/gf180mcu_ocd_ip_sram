magic
tech gf180mcuD
magscale 1 10
timestamp 1765480160
<< metal1 >>
rect -34 35 34 44
rect -34 -495 -26 35
rect 26 -495 34 35
rect -34 -504 34 -495
<< via1 >>
rect -26 -495 26 35
<< metal2 >>
rect -34 35 34 44
rect -34 -495 -26 35
rect 26 -495 34 35
rect -34 -504 34 -495
<< end >>
