magic
tech gf180mcuD
magscale 1 10
timestamp 1765484428
<< metal3 >>
rect -1397 77365 16227 77617
rect -1397 76651 16315 76903
rect -1397 76153 16315 76405
rect -1397 75439 16315 75691
rect -1397 74941 16315 75193
rect -1397 74227 16315 74479
rect -1397 73729 16315 73981
rect -1397 73015 16315 73267
rect -1397 72517 16315 72769
rect -1397 71803 16315 72055
rect -1397 71305 16315 71557
rect -1397 70591 16315 70843
rect -1397 70093 16315 70345
rect -1397 69379 16315 69631
rect -1397 68881 16315 69133
rect -1397 68167 16315 68419
rect -1397 67669 16315 67921
rect -1397 66955 16315 67207
rect -1397 66457 16315 66709
rect -1397 65743 16315 65995
rect -1397 65245 16315 65497
rect -1397 64531 16315 64783
rect -1397 64033 16315 64285
rect -1397 63319 16315 63571
rect -1397 62821 16315 63073
rect -1397 62107 16315 62359
rect -1397 61609 16315 61861
rect -1397 60895 16315 61147
rect -1397 60397 16315 60649
rect -1397 59683 16315 59935
rect -1397 59185 16315 59437
rect -1397 58471 16315 58723
rect -1397 57973 16315 58225
rect -1397 57259 16315 57511
rect -1397 56761 16315 57013
rect -1397 56047 16315 56299
rect -1397 55549 16315 55801
rect -1397 54835 16315 55087
rect -1397 54337 16315 54589
rect -1397 53623 16315 53875
rect -1397 53125 16315 53377
rect -1397 52411 16315 52663
rect -1397 51913 16315 52165
rect -1397 51199 16315 51451
rect -1397 50701 16315 50953
rect -1397 49987 16315 50239
rect -1397 49489 16315 49741
rect -1397 48775 16315 49027
rect -1397 48277 16315 48529
rect -1397 47563 16315 47815
rect -1397 47065 16315 47317
rect -1397 46351 16315 46603
rect -1397 45853 16315 46105
rect -1397 45139 16315 45391
rect -1397 44641 16315 44893
rect -1397 43927 16315 44179
rect -1397 43429 16315 43681
rect -1397 42715 16315 42967
rect -1397 42217 16315 42469
rect -1397 41503 16315 41755
rect -1397 41005 16315 41257
rect -1397 40291 16315 40543
rect -1397 39793 16315 40045
rect -1397 39079 16315 39331
rect -1397 38581 16315 38833
rect -1397 37867 16315 38119
rect -1397 37369 16315 37621
rect -1397 36906 -26 36907
rect 124 36906 16315 36907
rect -1397 36655 16315 36906
rect -26 36654 124 36655
rect -1397 36408 -26 36409
rect 124 36408 16315 36409
rect -1397 36157 16315 36408
rect -26 36156 124 36157
rect -1397 35694 -26 35695
rect 124 35694 16315 35695
rect -1397 35443 16315 35694
rect -26 35442 124 35443
rect -1397 35196 -26 35197
rect 124 35196 16315 35197
rect -1397 34945 16315 35196
rect -26 34944 124 34945
rect -1397 34482 -26 34483
rect 124 34482 16315 34483
rect -1397 34231 16315 34482
rect -26 34230 124 34231
rect -1397 33984 -26 33985
rect 124 33984 16315 33985
rect -1397 33733 16315 33984
rect -26 33732 124 33733
rect -1397 33270 -26 33271
rect 124 33270 16315 33271
rect -1397 33019 16315 33270
rect -26 33018 124 33019
rect -1397 32772 -26 32773
rect 124 32772 16315 32773
rect -1397 32521 16315 32772
rect -26 32520 124 32521
rect -1397 32058 -26 32059
rect 124 32058 16315 32059
rect -1397 31807 16315 32058
rect -26 31806 124 31807
rect -1397 31560 -26 31561
rect 124 31560 16315 31561
rect -1397 31309 16315 31560
rect -26 31308 124 31309
rect -1397 30846 -26 30847
rect 124 30846 16315 30847
rect -1397 30595 16315 30846
rect -26 30594 124 30595
rect -1397 30348 -26 30349
rect 124 30348 16315 30349
rect -1397 30097 16315 30348
rect -26 30096 124 30097
rect -1397 29634 -26 29635
rect 124 29634 16315 29635
rect -1397 29383 16315 29634
rect -26 29382 124 29383
rect -1397 29136 -26 29137
rect 124 29136 16315 29137
rect -1397 28885 16315 29136
rect -26 28884 124 28885
rect -1397 28422 -26 28423
rect 124 28422 16315 28423
rect -1397 28171 16315 28422
rect -26 28170 124 28171
rect -1397 27924 -26 27925
rect 124 27924 16315 27925
rect -1397 27673 16315 27924
rect -26 27672 124 27673
rect -1397 27210 -26 27211
rect 124 27210 16315 27211
rect -1397 26959 16315 27210
rect -26 26958 124 26959
rect -1397 26712 -26 26713
rect 124 26712 16315 26713
rect -1397 26461 16315 26712
rect -26 26460 124 26461
rect -1397 25998 -26 25999
rect 124 25998 16315 25999
rect -1397 25747 16315 25998
rect -26 25746 124 25747
rect -1397 25500 -26 25501
rect 124 25500 16315 25501
rect -1397 25249 16315 25500
rect -26 25248 124 25249
rect -1397 24786 -26 24787
rect 124 24786 16315 24787
rect -1397 24535 16315 24786
rect -26 24534 124 24535
rect -1397 24288 -26 24289
rect 124 24288 16315 24289
rect -1397 24037 16315 24288
rect -26 24036 124 24037
rect -1397 23574 -26 23575
rect 124 23574 16315 23575
rect -1397 23323 16315 23574
rect -26 23322 124 23323
rect -1397 23076 -26 23077
rect 124 23076 16315 23077
rect -1397 22825 16315 23076
rect -26 22824 124 22825
rect -1397 22362 -26 22363
rect 124 22362 16315 22363
rect -1397 22111 16315 22362
rect -26 22110 124 22111
rect -1397 21864 -26 21865
rect 124 21864 16315 21865
rect -1397 21613 16315 21864
rect -26 21612 124 21613
rect -1397 21150 -26 21151
rect 124 21150 16315 21151
rect -1397 20899 16315 21150
rect -26 20898 124 20899
rect -1397 20652 -26 20653
rect 124 20652 16315 20653
rect -1397 20401 16315 20652
rect -26 20400 124 20401
rect -1397 19938 -26 19939
rect 124 19938 16315 19939
rect -1397 19687 16315 19938
rect -26 19686 124 19687
rect -1397 19440 -26 19441
rect 124 19440 16315 19441
rect -1397 19189 16315 19440
rect -26 19188 124 19189
rect -1397 18726 -26 18727
rect 124 18726 16315 18727
rect -1397 18475 16315 18726
rect -26 18474 124 18475
rect -1397 18228 -26 18229
rect 124 18228 16315 18229
rect -1397 17977 16315 18228
rect -26 17976 124 17977
rect -1397 17514 -26 17515
rect 124 17514 16315 17515
rect -1397 17263 16315 17514
rect -26 17262 124 17263
rect -1397 17016 -26 17017
rect 124 17016 16315 17017
rect -1397 16765 16315 17016
rect -26 16764 124 16765
rect -1397 16302 -26 16303
rect 124 16302 16315 16303
rect -1397 16051 16315 16302
rect -26 16050 124 16051
rect -1397 15804 -26 15805
rect 124 15804 16315 15805
rect -1397 15553 16315 15804
rect -26 15552 124 15553
rect -1397 15090 -26 15091
rect 124 15090 16315 15091
rect -1397 14839 16315 15090
rect -26 14838 124 14839
rect -1397 14592 -26 14593
rect 124 14592 16315 14593
rect -1397 14341 16315 14592
rect -26 14340 124 14341
rect -1397 13878 -26 13879
rect 124 13878 16315 13879
rect -1397 13627 16315 13878
rect -26 13626 124 13627
rect -1397 13380 -26 13381
rect 124 13380 16315 13381
rect -1397 13129 16315 13380
rect -26 13128 124 13129
rect -1397 12666 -26 12667
rect 124 12666 16315 12667
rect -1397 12415 16315 12666
rect -26 12414 124 12415
rect -1397 12168 -26 12169
rect 124 12168 16315 12169
rect -1397 11917 16315 12168
rect -26 11916 124 11917
rect -1397 11454 -26 11455
rect 124 11454 16315 11455
rect -1397 11203 16315 11454
rect -26 11202 124 11203
rect -1397 10956 -26 10957
rect 124 10956 16315 10957
rect -1397 10705 16315 10956
rect -26 10704 124 10705
rect -1397 10242 -26 10243
rect 124 10242 16315 10243
rect -1397 9991 16315 10242
rect -26 9990 124 9991
rect -1397 9744 -26 9745
rect 124 9744 16315 9745
rect -1397 9493 16315 9744
rect -26 9492 124 9493
rect -1397 9030 -26 9031
rect 124 9030 16315 9031
rect -1397 8779 16315 9030
rect -26 8778 124 8779
rect -1397 8532 -26 8533
rect 124 8532 16315 8533
rect -1397 8281 16315 8532
rect -26 8280 124 8281
rect -1397 7818 -26 7819
rect 124 7818 16315 7819
rect -1397 7567 16315 7818
rect -26 7566 124 7567
rect -1397 7320 -26 7321
rect 124 7320 16315 7321
rect -1397 7069 16315 7320
rect -26 7068 124 7069
rect -1397 6606 -26 6607
rect 124 6606 16315 6607
rect -1397 6355 16315 6606
rect -26 6354 124 6355
rect -1397 6108 -26 6109
rect 124 6108 16315 6109
rect -1397 5857 16315 6108
rect -26 5856 124 5857
rect -1397 5394 -26 5395
rect 124 5394 16315 5395
rect -1397 5143 16315 5394
rect -26 5142 124 5143
rect -1397 4896 -26 4897
rect 124 4896 16315 4897
rect -1397 4645 16315 4896
rect -26 4644 124 4645
rect -1397 4182 -26 4183
rect 124 4182 16315 4183
rect -1397 3931 16315 4182
rect -26 3930 124 3931
rect -1397 3684 -26 3685
rect 124 3684 16315 3685
rect -1397 3433 16315 3684
rect -26 3432 124 3433
rect -1397 2970 -26 2971
rect 124 2970 16315 2971
rect -1397 2719 16315 2970
rect -26 2718 124 2719
rect -1397 2472 -26 2473
rect 124 2472 16315 2473
rect -1397 2221 16315 2472
rect -26 2220 124 2221
rect -1397 1758 -26 1759
rect 124 1758 16315 1759
rect -1397 1507 16315 1758
rect -26 1506 124 1507
rect -1397 1260 -26 1261
rect 124 1260 16315 1261
rect -1397 1009 16315 1260
rect -26 1008 124 1009
rect -1397 247 16315 499
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_0
timestamp 1764626446
transform -1 0 13007 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1
timestamp 1764626446
transform -1 0 13007 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2
timestamp 1764626446
transform -1 0 13007 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_3
timestamp 1764626446
transform -1 0 12571 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_4
timestamp 1764626446
transform -1 0 12571 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_5
timestamp 1764626446
transform -1 0 12571 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_6
timestamp 1764626446
transform -1 0 13007 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_7
timestamp 1764626446
transform -1 0 12571 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_8
timestamp 1764626446
transform -1 0 15623 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_9
timestamp 1764626446
transform -1 0 12571 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_10
timestamp 1764626446
transform -1 0 15623 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_11
timestamp 1764626446
transform -1 0 15623 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_12
timestamp 1764626446
transform -1 0 15623 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_13
timestamp 1764626446
transform -1 0 15623 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_14
timestamp 1764626446
transform -1 0 15623 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_15
timestamp 1764626446
transform -1 0 15623 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_16
timestamp 1764626446
transform -1 0 13443 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_17
timestamp 1764626446
transform -1 0 13879 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_18
timestamp 1764626446
transform -1 0 13879 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_19
timestamp 1764626446
transform -1 0 13879 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_20
timestamp 1764626446
transform -1 0 13879 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_21
timestamp 1764626446
transform -1 0 13879 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_22
timestamp 1764626446
transform -1 0 13879 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_23
timestamp 1764626446
transform -1 0 13879 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_24
timestamp 1764626446
transform -1 0 13443 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_25
timestamp 1764626446
transform -1 0 13007 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_26
timestamp 1764626446
transform -1 0 13443 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_27
timestamp 1764626446
transform -1 0 13007 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_28
timestamp 1764626446
transform -1 0 13443 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_29
timestamp 1764626446
transform -1 0 13443 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_30
timestamp 1764626446
transform -1 0 12571 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_31
timestamp 1764626446
transform -1 0 12571 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_32
timestamp 1764626446
transform -1 0 13443 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_33
timestamp 1764626446
transform -1 0 13443 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_34
timestamp 1764626446
transform -1 0 14751 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_35
timestamp 1764626446
transform -1 0 14751 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_36
timestamp 1764626446
transform -1 0 14315 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_37
timestamp 1764626446
transform -1 0 14315 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_38
timestamp 1764626446
transform -1 0 14315 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_39
timestamp 1764626446
transform -1 0 14315 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_40
timestamp 1764626446
transform -1 0 15187 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_41
timestamp 1764626446
transform -1 0 15187 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_42
timestamp 1764626446
transform -1 0 15187 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_43
timestamp 1764626446
transform -1 0 15187 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_44
timestamp 1764626446
transform -1 0 15187 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_45
timestamp 1764626446
transform -1 0 15187 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_46
timestamp 1764626446
transform -1 0 15187 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_47
timestamp 1764626446
transform -1 0 14315 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_48
timestamp 1764626446
transform -1 0 14315 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_49
timestamp 1764626446
transform -1 0 14315 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_50
timestamp 1764626446
transform -1 0 13007 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_51
timestamp 1764626446
transform -1 0 14751 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_52
timestamp 1764626446
transform -1 0 14751 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_53
timestamp 1764626446
transform -1 0 14751 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_54
timestamp 1764626446
transform -1 0 14751 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_55
timestamp 1764626446
transform -1 0 14751 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_56
timestamp 1764626446
transform 1 0 8063 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_57
timestamp 1764626446
transform 1 0 8063 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_58
timestamp 1764626446
transform 1 0 8063 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_59
timestamp 1764626446
transform 1 0 8063 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_60
timestamp 1764626446
transform 1 0 8063 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_61
timestamp 1764626446
transform 1 0 8063 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_62
timestamp 1764626446
transform 1 0 8063 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_63
timestamp 1764626446
transform 1 0 8499 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_64
timestamp 1764626446
transform 1 0 8499 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_65
timestamp 1764626446
transform 1 0 8499 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_66
timestamp 1764626446
transform 1 0 10679 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_67
timestamp 1764626446
transform 1 0 10243 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_68
timestamp 1764626446
transform 1 0 10679 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_69
timestamp 1764626446
transform 1 0 10679 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_70
timestamp 1764626446
transform 1 0 10679 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_71
timestamp 1764626446
transform 1 0 10679 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_72
timestamp 1764626446
transform 1 0 8935 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_73
timestamp 1764626446
transform 1 0 8935 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_74
timestamp 1764626446
transform 1 0 8935 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_75
timestamp 1764626446
transform 1 0 8935 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_76
timestamp 1764626446
transform 1 0 10243 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_77
timestamp 1764626446
transform 1 0 10243 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_78
timestamp 1764626446
transform 1 0 10243 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_79
timestamp 1764626446
transform 1 0 10243 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_80
timestamp 1764626446
transform 1 0 10243 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_81
timestamp 1764626446
transform 1 0 10243 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_82
timestamp 1764626446
transform 1 0 8935 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_83
timestamp 1764626446
transform 1 0 10679 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_84
timestamp 1764626446
transform 1 0 9807 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_85
timestamp 1764626446
transform 1 0 9807 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_86
timestamp 1764626446
transform 1 0 9807 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_87
timestamp 1764626446
transform 1 0 9807 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_88
timestamp 1764626446
transform 1 0 9807 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_89
timestamp 1764626446
transform 1 0 10679 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_90
timestamp 1764626446
transform 1 0 11115 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_91
timestamp 1764626446
transform 1 0 11115 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_92
timestamp 1764626446
transform 1 0 11115 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_93
timestamp 1764626446
transform 1 0 11115 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_94
timestamp 1764626446
transform 1 0 11115 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_95
timestamp 1764626446
transform 1 0 11115 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_96
timestamp 1764626446
transform 1 0 11115 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_97
timestamp 1764626446
transform 1 0 9807 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_98
timestamp 1764626446
transform 1 0 9807 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_99
timestamp 1764626446
transform 1 0 9371 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_100
timestamp 1764626446
transform 1 0 9371 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_101
timestamp 1764626446
transform 1 0 9371 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_102
timestamp 1764626446
transform 1 0 9371 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_103
timestamp 1764626446
transform 1 0 9371 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_104
timestamp 1764626446
transform 1 0 9371 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_105
timestamp 1764626446
transform 1 0 9371 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_106
timestamp 1764626446
transform 1 0 8499 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_107
timestamp 1764626446
transform 1 0 8499 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_108
timestamp 1764626446
transform 1 0 8499 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_109
timestamp 1764626446
transform 1 0 8499 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_110
timestamp 1764626446
transform 1 0 8935 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_111
timestamp 1764626446
transform 1 0 8935 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_112
timestamp 1764626446
transform 1 0 11115 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_113
timestamp 1764626446
transform 1 0 8063 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_114
timestamp 1764626446
transform 1 0 11115 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_115
timestamp 1764626446
transform 1 0 11115 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_116
timestamp 1764626446
transform 1 0 11115 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_117
timestamp 1764626446
transform 1 0 9371 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_118
timestamp 1764626446
transform 1 0 11115 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_119
timestamp 1764626446
transform 1 0 9371 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_120
timestamp 1764626446
transform 1 0 8063 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_121
timestamp 1764626446
transform 1 0 8063 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_122
timestamp 1764626446
transform 1 0 9371 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_123
timestamp 1764626446
transform 1 0 10679 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_124
timestamp 1764626446
transform 1 0 10679 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_125
timestamp 1764626446
transform 1 0 9371 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_126
timestamp 1764626446
transform 1 0 9371 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_127
timestamp 1764626446
transform 1 0 8499 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_128
timestamp 1764626446
transform 1 0 8499 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_129
timestamp 1764626446
transform 1 0 10679 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_130
timestamp 1764626446
transform 1 0 10679 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_131
timestamp 1764626446
transform 1 0 10679 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_132
timestamp 1764626446
transform 1 0 10679 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_133
timestamp 1764626446
transform 1 0 9371 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_134
timestamp 1764626446
transform 1 0 11115 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_135
timestamp 1764626446
transform 1 0 8499 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_136
timestamp 1764626446
transform 1 0 8935 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_137
timestamp 1764626446
transform 1 0 10243 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_138
timestamp 1764626446
transform 1 0 10243 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_139
timestamp 1764626446
transform 1 0 10243 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_140
timestamp 1764626446
transform 1 0 10243 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_141
timestamp 1764626446
transform 1 0 10243 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_142
timestamp 1764626446
transform 1 0 10243 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_143
timestamp 1764626446
transform 1 0 8063 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_144
timestamp 1764626446
transform 1 0 8063 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_145
timestamp 1764626446
transform 1 0 8935 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_146
timestamp 1764626446
transform 1 0 8935 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_147
timestamp 1764626446
transform 1 0 8935 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_148
timestamp 1764626446
transform 1 0 8935 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_149
timestamp 1764626446
transform 1 0 8935 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_150
timestamp 1764626446
transform 1 0 9807 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_151
timestamp 1764626446
transform 1 0 9807 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_152
timestamp 1764626446
transform 1 0 9807 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_153
timestamp 1764626446
transform 1 0 9807 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_154
timestamp 1764626446
transform 1 0 9807 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_155
timestamp 1764626446
transform 1 0 9807 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_156
timestamp 1764626446
transform 1 0 8499 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_157
timestamp 1764626446
transform 1 0 8499 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_158
timestamp 1764626446
transform 1 0 8499 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_159
timestamp 1764626446
transform 1 0 8063 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_160
timestamp 1764626446
transform -1 0 13007 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_161
timestamp 1764626446
transform -1 0 14751 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_162
timestamp 1764626446
transform -1 0 13007 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_163
timestamp 1764626446
transform -1 0 13007 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_164
timestamp 1764626446
transform -1 0 13007 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_165
timestamp 1764626446
transform -1 0 13007 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_166
timestamp 1764626446
transform -1 0 13007 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_167
timestamp 1764626446
transform -1 0 14751 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_168
timestamp 1764626446
transform -1 0 14315 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_169
timestamp 1764626446
transform -1 0 14315 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_170
timestamp 1764626446
transform -1 0 13443 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_171
timestamp 1764626446
transform -1 0 12571 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_172
timestamp 1764626446
transform -1 0 12571 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_173
timestamp 1764626446
transform -1 0 12571 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_174
timestamp 1764626446
transform -1 0 12571 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_175
timestamp 1764626446
transform -1 0 12571 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_176
timestamp 1764626446
transform -1 0 12571 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_177
timestamp 1764626446
transform -1 0 13443 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_178
timestamp 1764626446
transform -1 0 13443 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_179
timestamp 1764626446
transform -1 0 13443 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_180
timestamp 1764626446
transform -1 0 13443 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_181
timestamp 1764626446
transform -1 0 13443 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_182
timestamp 1764626446
transform -1 0 14315 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_183
timestamp 1764626446
transform -1 0 15623 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_184
timestamp 1764626446
transform -1 0 15623 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_185
timestamp 1764626446
transform -1 0 15623 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_186
timestamp 1764626446
transform -1 0 15623 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_187
timestamp 1764626446
transform -1 0 15623 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_188
timestamp 1764626446
transform -1 0 15623 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_189
timestamp 1764626446
transform -1 0 14315 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_190
timestamp 1764626446
transform -1 0 14315 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_191
timestamp 1764626446
transform -1 0 14315 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_192
timestamp 1764626446
transform -1 0 14751 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_193
timestamp 1764626446
transform -1 0 15187 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_194
timestamp 1764626446
transform -1 0 15187 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_195
timestamp 1764626446
transform -1 0 15187 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_196
timestamp 1764626446
transform -1 0 15187 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_197
timestamp 1764626446
transform -1 0 15187 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_198
timestamp 1764626446
transform -1 0 15187 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_199
timestamp 1764626446
transform -1 0 14751 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_200
timestamp 1764626446
transform -1 0 14751 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_201
timestamp 1764626446
transform -1 0 14751 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_202
timestamp 1764626446
transform -1 0 13879 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_203
timestamp 1764626446
transform -1 0 13879 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_204
timestamp 1764626446
transform -1 0 13879 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_205
timestamp 1764626446
transform -1 0 13879 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_206
timestamp 1764626446
transform -1 0 13879 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_207
timestamp 1764626446
transform -1 0 13879 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_208
timestamp 1764626446
transform -1 0 13007 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_209
timestamp 1764626446
transform -1 0 13007 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_210
timestamp 1764626446
transform -1 0 12571 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_211
timestamp 1764626446
transform -1 0 12571 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_212
timestamp 1764626446
transform 1 0 9807 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_213
timestamp 1764626446
transform 1 0 9807 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_214
timestamp 1764626446
transform 1 0 8063 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_215
timestamp 1764626446
transform 1 0 8063 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_216
timestamp 1764626446
transform -1 0 15623 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_217
timestamp 1764626446
transform -1 0 15623 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_218
timestamp 1764626446
transform 1 0 10243 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_219
timestamp 1764626446
transform 1 0 10243 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_220
timestamp 1764626446
transform -1 0 15187 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_221
timestamp 1764626446
transform -1 0 15187 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_222
timestamp 1764626446
transform -1 0 13879 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_223
timestamp 1764626446
transform -1 0 13879 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_224
timestamp 1764626446
transform 1 0 8935 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_225
timestamp 1764626446
transform 1 0 8935 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_226
timestamp 1764626446
transform -1 0 13443 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_227
timestamp 1764626446
transform -1 0 13443 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_228
timestamp 1764626446
transform 1 0 10679 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_229
timestamp 1764626446
transform 1 0 10679 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_230
timestamp 1764626446
transform -1 0 14751 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_231
timestamp 1764626446
transform -1 0 14751 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_232
timestamp 1764626446
transform 1 0 8499 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_233
timestamp 1764626446
transform 1 0 8499 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_234
timestamp 1764626446
transform -1 0 14315 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_235
timestamp 1764626446
transform -1 0 14315 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_236
timestamp 1764626446
transform 1 0 9371 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_237
timestamp 1764626446
transform 1 0 9371 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_238
timestamp 1764626446
transform 1 0 11115 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_239
timestamp 1764626446
transform 1 0 11115 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_240
timestamp 1764626446
transform -1 0 6935 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_241
timestamp 1764626446
transform -1 0 6935 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_242
timestamp 1764626446
transform -1 0 6935 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_243
timestamp 1764626446
transform -1 0 6935 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_244
timestamp 1764626446
transform -1 0 6935 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_245
timestamp 1764626446
transform -1 0 6935 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_246
timestamp 1764626446
transform -1 0 6935 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_247
timestamp 1764626446
transform -1 0 7807 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_248
timestamp 1764626446
transform -1 0 7807 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_249
timestamp 1764626446
transform -1 0 7807 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_250
timestamp 1764626446
transform -1 0 5627 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_251
timestamp 1764626446
transform -1 0 5627 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_252
timestamp 1764626446
transform -1 0 5627 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_253
timestamp 1764626446
transform -1 0 5627 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_254
timestamp 1764626446
transform -1 0 5627 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_255
timestamp 1764626446
transform -1 0 5627 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_256
timestamp 1764626446
transform -1 0 5627 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_257
timestamp 1764626446
transform -1 0 4755 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_258
timestamp 1764626446
transform -1 0 4755 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_259
timestamp 1764626446
transform -1 0 4755 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_260
timestamp 1764626446
transform -1 0 4755 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_261
timestamp 1764626446
transform -1 0 4755 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_262
timestamp 1764626446
transform -1 0 4755 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_263
timestamp 1764626446
transform -1 0 4755 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_264
timestamp 1764626446
transform -1 0 7807 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_265
timestamp 1764626446
transform -1 0 7807 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_266
timestamp 1764626446
transform -1 0 7807 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_267
timestamp 1764626446
transform -1 0 7807 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_268
timestamp 1764626446
transform -1 0 7371 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_269
timestamp 1764626446
transform -1 0 7371 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_270
timestamp 1764626446
transform -1 0 7371 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_271
timestamp 1764626446
transform -1 0 7371 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_272
timestamp 1764626446
transform -1 0 7371 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_273
timestamp 1764626446
transform -1 0 7371 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_274
timestamp 1764626446
transform -1 0 7371 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_275
timestamp 1764626446
transform -1 0 6063 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_276
timestamp 1764626446
transform -1 0 6063 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_277
timestamp 1764626446
transform -1 0 6063 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_278
timestamp 1764626446
transform -1 0 6499 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_279
timestamp 1764626446
transform -1 0 6499 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_280
timestamp 1764626446
transform -1 0 6499 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_281
timestamp 1764626446
transform -1 0 6499 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_282
timestamp 1764626446
transform -1 0 5191 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_283
timestamp 1764626446
transform -1 0 5191 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_284
timestamp 1764626446
transform -1 0 5191 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_285
timestamp 1764626446
transform -1 0 5191 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_286
timestamp 1764626446
transform -1 0 5191 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_287
timestamp 1764626446
transform -1 0 5191 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_288
timestamp 1764626446
transform -1 0 5191 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_289
timestamp 1764626446
transform -1 0 6499 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_290
timestamp 1764626446
transform -1 0 6499 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_291
timestamp 1764626446
transform -1 0 6499 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_292
timestamp 1764626446
transform -1 0 6063 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_293
timestamp 1764626446
transform -1 0 6063 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_294
timestamp 1764626446
transform -1 0 6063 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_295
timestamp 1764626446
transform -1 0 6063 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_296
timestamp 1764626446
transform 1 0 1119 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_297
timestamp 1764626446
transform 1 0 247 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_298
timestamp 1764626446
transform 1 0 247 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_299
timestamp 1764626446
transform 1 0 247 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_300
timestamp 1764626446
transform 1 0 1555 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_301
timestamp 1764626446
transform 1 0 1555 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_302
timestamp 1764626446
transform 1 0 1555 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_303
timestamp 1764626446
transform 1 0 1555 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_304
timestamp 1764626446
transform 1 0 1555 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_305
timestamp 1764626446
transform 1 0 1555 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_306
timestamp 1764626446
transform 1 0 247 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_307
timestamp 1764626446
transform 1 0 247 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_308
timestamp 1764626446
transform 1 0 247 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_309
timestamp 1764626446
transform 1 0 683 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_310
timestamp 1764626446
transform 1 0 683 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_311
timestamp 1764626446
transform 1 0 683 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_312
timestamp 1764626446
transform 1 0 3299 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_313
timestamp 1764626446
transform 1 0 3299 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_314
timestamp 1764626446
transform 1 0 3299 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_315
timestamp 1764626446
transform 1 0 3299 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_316
timestamp 1764626446
transform 1 0 3299 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_317
timestamp 1764626446
transform 1 0 3299 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_318
timestamp 1764626446
transform 1 0 3299 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_319
timestamp 1764626446
transform 1 0 683 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_320
timestamp 1764626446
transform 1 0 683 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_321
timestamp 1764626446
transform 1 0 2863 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_322
timestamp 1764626446
transform 1 0 2863 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_323
timestamp 1764626446
transform 1 0 2863 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_324
timestamp 1764626446
transform 1 0 2863 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_325
timestamp 1764626446
transform 1 0 2863 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_326
timestamp 1764626446
transform 1 0 683 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_327
timestamp 1764626446
transform 1 0 1991 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_328
timestamp 1764626446
transform 1 0 1991 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_329
timestamp 1764626446
transform 1 0 1991 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_330
timestamp 1764626446
transform 1 0 1991 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_331
timestamp 1764626446
transform 1 0 2863 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_332
timestamp 1764626446
transform 1 0 2863 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_333
timestamp 1764626446
transform 1 0 1991 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_334
timestamp 1764626446
transform 1 0 1991 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_335
timestamp 1764626446
transform 1 0 1991 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_336
timestamp 1764626446
transform 1 0 2427 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_337
timestamp 1764626446
transform 1 0 2427 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_338
timestamp 1764626446
transform 1 0 2427 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_339
timestamp 1764626446
transform 1 0 2427 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_340
timestamp 1764626446
transform 1 0 2427 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_341
timestamp 1764626446
transform 1 0 1555 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_342
timestamp 1764626446
transform 1 0 2427 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_343
timestamp 1764626446
transform 1 0 2427 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_344
timestamp 1764626446
transform 1 0 683 0 1 7272
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_345
timestamp 1764626446
transform 1 0 1119 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_346
timestamp 1764626446
transform 1 0 247 0 1 1212
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_347
timestamp 1764626446
transform 1 0 1119 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_348
timestamp 1764626446
transform 1 0 1119 0 1 2424
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_349
timestamp 1764626446
transform 1 0 1119 0 1 3636
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_350
timestamp 1764626446
transform 1 0 1119 0 1 4848
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_351
timestamp 1764626446
transform 1 0 1119 0 1 6060
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_352
timestamp 1764626446
transform 1 0 683 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_353
timestamp 1764626446
transform 1 0 683 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_354
timestamp 1764626446
transform 1 0 683 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_355
timestamp 1764626446
transform 1 0 3299 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_356
timestamp 1764626446
transform 1 0 3299 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_357
timestamp 1764626446
transform 1 0 3299 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_358
timestamp 1764626446
transform 1 0 3299 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_359
timestamp 1764626446
transform 1 0 3299 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_360
timestamp 1764626446
transform 1 0 1555 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_361
timestamp 1764626446
transform 1 0 1555 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_362
timestamp 1764626446
transform 1 0 1555 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_363
timestamp 1764626446
transform 1 0 1555 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_364
timestamp 1764626446
transform 1 0 1555 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_365
timestamp 1764626446
transform 1 0 1555 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_366
timestamp 1764626446
transform 1 0 2427 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_367
timestamp 1764626446
transform 1 0 2427 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_368
timestamp 1764626446
transform 1 0 2427 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_369
timestamp 1764626446
transform 1 0 2427 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_370
timestamp 1764626446
transform 1 0 2427 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_371
timestamp 1764626446
transform 1 0 683 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_372
timestamp 1764626446
transform 1 0 683 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_373
timestamp 1764626446
transform 1 0 3299 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_374
timestamp 1764626446
transform 1 0 247 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_375
timestamp 1764626446
transform 1 0 247 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_376
timestamp 1764626446
transform 1 0 247 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_377
timestamp 1764626446
transform 1 0 247 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_378
timestamp 1764626446
transform 1 0 2427 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_379
timestamp 1764626446
transform 1 0 1119 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_380
timestamp 1764626446
transform 1 0 2863 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_381
timestamp 1764626446
transform 1 0 2863 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_382
timestamp 1764626446
transform 1 0 2863 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_383
timestamp 1764626446
transform 1 0 2863 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_384
timestamp 1764626446
transform 1 0 2863 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_385
timestamp 1764626446
transform 1 0 2863 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_386
timestamp 1764626446
transform 1 0 1991 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_387
timestamp 1764626446
transform 1 0 1991 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_388
timestamp 1764626446
transform 1 0 1991 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_389
timestamp 1764626446
transform 1 0 1991 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_390
timestamp 1764626446
transform 1 0 1991 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_391
timestamp 1764626446
transform 1 0 1991 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_392
timestamp 1764626446
transform 1 0 247 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_393
timestamp 1764626446
transform 1 0 247 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_394
timestamp 1764626446
transform 1 0 1119 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_395
timestamp 1764626446
transform 1 0 1119 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_396
timestamp 1764626446
transform 1 0 1119 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_397
timestamp 1764626446
transform 1 0 1119 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_398
timestamp 1764626446
transform 1 0 1119 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_399
timestamp 1764626446
transform 1 0 683 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_400
timestamp 1764626446
transform -1 0 7371 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_401
timestamp 1764626446
transform -1 0 7371 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_402
timestamp 1764626446
transform -1 0 7371 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_403
timestamp 1764626446
transform -1 0 7371 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_404
timestamp 1764626446
transform -1 0 7371 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_405
timestamp 1764626446
transform -1 0 7371 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_406
timestamp 1764626446
transform -1 0 7807 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_407
timestamp 1764626446
transform -1 0 7807 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_408
timestamp 1764626446
transform -1 0 7807 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_409
timestamp 1764626446
transform -1 0 6063 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_410
timestamp 1764626446
transform -1 0 6063 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_411
timestamp 1764626446
transform -1 0 5191 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_412
timestamp 1764626446
transform -1 0 5191 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_413
timestamp 1764626446
transform -1 0 5191 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_414
timestamp 1764626446
transform -1 0 5191 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_415
timestamp 1764626446
transform -1 0 5191 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_416
timestamp 1764626446
transform -1 0 5191 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_417
timestamp 1764626446
transform -1 0 6063 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_418
timestamp 1764626446
transform -1 0 6063 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_419
timestamp 1764626446
transform -1 0 6063 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_420
timestamp 1764626446
transform -1 0 6063 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_421
timestamp 1764626446
transform -1 0 4755 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_422
timestamp 1764626446
transform -1 0 4755 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_423
timestamp 1764626446
transform -1 0 4755 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_424
timestamp 1764626446
transform -1 0 4755 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_425
timestamp 1764626446
transform -1 0 4755 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_426
timestamp 1764626446
transform -1 0 4755 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_427
timestamp 1764626446
transform -1 0 7807 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_428
timestamp 1764626446
transform -1 0 7807 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_429
timestamp 1764626446
transform -1 0 7807 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_430
timestamp 1764626446
transform -1 0 5627 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_431
timestamp 1764626446
transform -1 0 6935 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_432
timestamp 1764626446
transform -1 0 6935 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_433
timestamp 1764626446
transform -1 0 6935 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_434
timestamp 1764626446
transform -1 0 6935 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_435
timestamp 1764626446
transform -1 0 6935 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_436
timestamp 1764626446
transform -1 0 6935 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_437
timestamp 1764626446
transform -1 0 5627 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_438
timestamp 1764626446
transform -1 0 5627 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_439
timestamp 1764626446
transform -1 0 5627 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_440
timestamp 1764626446
transform -1 0 5627 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_441
timestamp 1764626446
transform -1 0 6499 0 1 10908
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_442
timestamp 1764626446
transform -1 0 6499 0 1 12120
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_443
timestamp 1764626446
transform -1 0 6499 0 1 13332
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_444
timestamp 1764626446
transform -1 0 6499 0 1 14544
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_445
timestamp 1764626446
transform -1 0 6499 0 1 15756
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_446
timestamp 1764626446
transform -1 0 6499 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_447
timestamp 1764626446
transform -1 0 5627 0 1 16968
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_448
timestamp 1764626446
transform 1 0 1555 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_449
timestamp 1764626446
transform 1 0 1555 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_450
timestamp 1764626446
transform -1 0 5191 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_451
timestamp 1764626446
transform -1 0 5191 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_452
timestamp 1764626446
transform 1 0 2863 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_453
timestamp 1764626446
transform 1 0 2863 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_454
timestamp 1764626446
transform -1 0 4755 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_455
timestamp 1764626446
transform -1 0 4755 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_456
timestamp 1764626446
transform 1 0 247 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_457
timestamp 1764626446
transform 1 0 247 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_458
timestamp 1764626446
transform -1 0 6935 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_459
timestamp 1764626446
transform -1 0 6935 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_460
timestamp 1764626446
transform 1 0 3299 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_461
timestamp 1764626446
transform 1 0 3299 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_462
timestamp 1764626446
transform -1 0 6499 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_463
timestamp 1764626446
transform -1 0 6499 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_464
timestamp 1764626446
transform 1 0 1991 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_465
timestamp 1764626446
transform -1 0 6063 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_466
timestamp 1764626446
transform -1 0 6063 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_467
timestamp 1764626446
transform 1 0 1991 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_468
timestamp 1764626446
transform -1 0 5627 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_469
timestamp 1764626446
transform -1 0 5627 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_470
timestamp 1764626446
transform 1 0 1119 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_471
timestamp 1764626446
transform 1 0 1119 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_472
timestamp 1764626446
transform 1 0 683 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_473
timestamp 1764626446
transform -1 0 7807 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_474
timestamp 1764626446
transform -1 0 7807 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_475
timestamp 1764626446
transform 1 0 683 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_476
timestamp 1764626446
transform 1 0 2427 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_477
timestamp 1764626446
transform 1 0 2427 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_478
timestamp 1764626446
transform -1 0 7371 0 1 8484
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_479
timestamp 1764626446
transform -1 0 7371 0 1 9696
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_480
timestamp 1764626446
transform -1 0 5191 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_481
timestamp 1764626446
transform -1 0 6499 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_482
timestamp 1764626446
transform -1 0 5627 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_483
timestamp 1764626446
transform -1 0 7371 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_484
timestamp 1764626446
transform -1 0 6063 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_485
timestamp 1764626446
transform -1 0 7371 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_486
timestamp 1764626446
transform -1 0 7807 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_487
timestamp 1764626446
transform -1 0 7807 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_488
timestamp 1764626446
transform -1 0 7807 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_489
timestamp 1764626446
transform -1 0 7807 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_490
timestamp 1764626446
transform -1 0 6499 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_491
timestamp 1764626446
transform -1 0 6499 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_492
timestamp 1764626446
transform -1 0 6499 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_493
timestamp 1764626446
transform -1 0 6499 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_494
timestamp 1764626446
transform -1 0 6499 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_495
timestamp 1764626446
transform -1 0 4755 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_496
timestamp 1764626446
transform -1 0 4755 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_497
timestamp 1764626446
transform -1 0 4755 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_498
timestamp 1764626446
transform -1 0 4755 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_499
timestamp 1764626446
transform -1 0 4755 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_500
timestamp 1764626446
transform -1 0 4755 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_501
timestamp 1764626446
transform -1 0 7807 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_502
timestamp 1764626446
transform -1 0 7371 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_503
timestamp 1764626446
transform -1 0 7371 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_504
timestamp 1764626446
transform -1 0 7371 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_505
timestamp 1764626446
transform -1 0 7807 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_506
timestamp 1764626446
transform -1 0 7371 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_507
timestamp 1764626446
transform -1 0 5627 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_508
timestamp 1764626446
transform -1 0 5627 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_509
timestamp 1764626446
transform -1 0 5627 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_510
timestamp 1764626446
transform -1 0 6935 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_511
timestamp 1764626446
transform -1 0 6063 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_512
timestamp 1764626446
transform -1 0 15623 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_513
timestamp 1764626446
transform -1 0 6935 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_514
timestamp 1764626446
transform -1 0 6935 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_515
timestamp 1764626446
transform -1 0 6935 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_516
timestamp 1764626446
transform -1 0 6935 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_517
timestamp 1764626446
transform -1 0 6935 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_518
timestamp 1764626446
transform -1 0 5627 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_519
timestamp 1764626446
transform -1 0 6063 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_520
timestamp 1764626446
transform -1 0 6063 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_521
timestamp 1764626446
transform -1 0 5191 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_522
timestamp 1764626446
transform -1 0 6063 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_523
timestamp 1764626446
transform -1 0 6063 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_524
timestamp 1764626446
transform -1 0 5191 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_525
timestamp 1764626446
transform -1 0 5191 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_526
timestamp 1764626446
transform -1 0 5191 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_527
timestamp 1764626446
transform -1 0 5191 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_528
timestamp 1764626446
transform 1 0 3299 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_529
timestamp 1764626446
transform 1 0 2427 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_530
timestamp 1764626446
transform 1 0 683 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_531
timestamp 1764626446
transform 1 0 1119 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_532
timestamp 1764626446
transform 1 0 1119 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_533
timestamp 1764626446
transform 1 0 1119 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_534
timestamp 1764626446
transform 1 0 1119 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_535
timestamp 1764626446
transform 1 0 1119 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_536
timestamp 1764626446
transform 1 0 1119 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_537
timestamp 1764626446
transform 1 0 1991 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_538
timestamp 1764626446
transform 1 0 1555 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_539
timestamp 1764626446
transform 1 0 2863 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_540
timestamp 1764626446
transform 1 0 1555 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_541
timestamp 1764626446
transform 1 0 1555 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_542
timestamp 1764626446
transform 1 0 1555 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_543
timestamp 1764626446
transform 1 0 1555 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_544
timestamp 1764626446
transform 1 0 1555 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_545
timestamp 1764626446
transform 1 0 2863 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_546
timestamp 1764626446
transform 1 0 683 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_547
timestamp 1764626446
transform 1 0 1991 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_548
timestamp 1764626446
transform 1 0 1991 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_549
timestamp 1764626446
transform 1 0 1991 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_550
timestamp 1764626446
transform 1 0 1991 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_551
timestamp 1764626446
transform 1 0 1991 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_552
timestamp 1764626446
transform 1 0 247 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_553
timestamp 1764626446
transform 1 0 683 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_554
timestamp 1764626446
transform 1 0 2863 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_555
timestamp 1764626446
transform 1 0 683 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_556
timestamp 1764626446
transform 1 0 247 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_557
timestamp 1764626446
transform 1 0 247 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_558
timestamp 1764626446
transform 1 0 247 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_559
timestamp 1764626446
transform 1 0 247 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_560
timestamp 1764626446
transform 1 0 247 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_561
timestamp 1764626446
transform 1 0 683 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_562
timestamp 1764626446
transform 1 0 683 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_563
timestamp 1764626446
transform 1 0 2427 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_564
timestamp 1764626446
transform 1 0 2863 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_565
timestamp 1764626446
transform 1 0 2427 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_566
timestamp 1764626446
transform 1 0 2427 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_567
timestamp 1764626446
transform 1 0 3299 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_568
timestamp 1764626446
transform 1 0 3299 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_569
timestamp 1764626446
transform 1 0 3299 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_570
timestamp 1764626446
transform 1 0 3299 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_571
timestamp 1764626446
transform 1 0 3299 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_572
timestamp 1764626446
transform 1 0 2427 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_573
timestamp 1764626446
transform 1 0 2427 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_574
timestamp 1764626446
transform 1 0 2863 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_575
timestamp 1764626446
transform 1 0 2863 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_576
timestamp 1764626446
transform 1 0 2427 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_577
timestamp 1764626446
transform 1 0 2427 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_578
timestamp 1764626446
transform 1 0 1119 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_579
timestamp 1764626446
transform 1 0 1119 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_580
timestamp 1764626446
transform 1 0 1119 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_581
timestamp 1764626446
transform 1 0 1119 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_582
timestamp 1764626446
transform 1 0 1119 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_583
timestamp 1764626446
transform 1 0 1119 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_584
timestamp 1764626446
transform 1 0 1119 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_585
timestamp 1764626446
transform 1 0 2427 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_586
timestamp 1764626446
transform 1 0 2427 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_587
timestamp 1764626446
transform 1 0 1555 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_588
timestamp 1764626446
transform 1 0 1555 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_589
timestamp 1764626446
transform 1 0 1555 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_590
timestamp 1764626446
transform 1 0 1555 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_591
timestamp 1764626446
transform 1 0 1555 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_592
timestamp 1764626446
transform 1 0 1555 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_593
timestamp 1764626446
transform 1 0 1555 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_594
timestamp 1764626446
transform 1 0 2427 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_595
timestamp 1764626446
transform 1 0 2427 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_596
timestamp 1764626446
transform 1 0 2863 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_597
timestamp 1764626446
transform 1 0 2863 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_598
timestamp 1764626446
transform 1 0 2427 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_599
timestamp 1764626446
transform 1 0 247 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_600
timestamp 1764626446
transform 1 0 247 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_601
timestamp 1764626446
transform 1 0 247 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_602
timestamp 1764626446
transform 1 0 247 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_603
timestamp 1764626446
transform 1 0 2863 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_604
timestamp 1764626446
transform 1 0 2863 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_605
timestamp 1764626446
transform 1 0 247 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_606
timestamp 1764626446
transform 1 0 247 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_607
timestamp 1764626446
transform 1 0 247 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_608
timestamp 1764626446
transform 1 0 683 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_609
timestamp 1764626446
transform 1 0 683 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_610
timestamp 1764626446
transform 1 0 2863 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_611
timestamp 1764626446
transform 1 0 683 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_612
timestamp 1764626446
transform 1 0 683 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_613
timestamp 1764626446
transform 1 0 3299 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_614
timestamp 1764626446
transform 1 0 3299 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_615
timestamp 1764626446
transform 1 0 3299 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_616
timestamp 1764626446
transform 1 0 3299 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_617
timestamp 1764626446
transform 1 0 3299 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_618
timestamp 1764626446
transform 1 0 3299 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_619
timestamp 1764626446
transform 1 0 3299 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_620
timestamp 1764626446
transform 1 0 683 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_621
timestamp 1764626446
transform 1 0 683 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_622
timestamp 1764626446
transform 1 0 1991 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_623
timestamp 1764626446
transform 1 0 1991 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_624
timestamp 1764626446
transform 1 0 1991 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_625
timestamp 1764626446
transform 1 0 1991 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_626
timestamp 1764626446
transform 1 0 1991 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_627
timestamp 1764626446
transform 1 0 1991 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_628
timestamp 1764626446
transform 1 0 1991 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_629
timestamp 1764626446
transform 1 0 2863 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_630
timestamp 1764626446
transform 1 0 2863 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_631
timestamp 1764626446
transform 1 0 683 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_632
timestamp 1764626446
transform -1 0 5627 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_633
timestamp 1764626446
transform -1 0 5627 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_634
timestamp 1764626446
transform -1 0 5627 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_635
timestamp 1764626446
transform -1 0 5627 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_636
timestamp 1764626446
transform -1 0 5627 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_637
timestamp 1764626446
transform -1 0 7371 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_638
timestamp 1764626446
transform -1 0 5191 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_639
timestamp 1764626446
transform -1 0 5191 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_640
timestamp 1764626446
transform -1 0 5191 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_641
timestamp 1764626446
transform -1 0 5191 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_642
timestamp 1764626446
transform -1 0 5191 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_643
timestamp 1764626446
transform -1 0 5191 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_644
timestamp 1764626446
transform -1 0 5191 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_645
timestamp 1764626446
transform -1 0 7371 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_646
timestamp 1764626446
transform -1 0 7807 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_647
timestamp 1764626446
transform -1 0 7807 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_648
timestamp 1764626446
transform -1 0 4755 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_649
timestamp 1764626446
transform -1 0 4755 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_650
timestamp 1764626446
transform -1 0 4755 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_651
timestamp 1764626446
transform -1 0 4755 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_652
timestamp 1764626446
transform -1 0 4755 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_653
timestamp 1764626446
transform -1 0 4755 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_654
timestamp 1764626446
transform -1 0 4755 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_655
timestamp 1764626446
transform -1 0 7807 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_656
timestamp 1764626446
transform -1 0 7807 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_657
timestamp 1764626446
transform -1 0 6935 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_658
timestamp 1764626446
transform -1 0 6935 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_659
timestamp 1764626446
transform -1 0 6935 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_660
timestamp 1764626446
transform -1 0 6935 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_661
timestamp 1764626446
transform -1 0 6935 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_662
timestamp 1764626446
transform -1 0 6935 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_663
timestamp 1764626446
transform -1 0 6935 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_664
timestamp 1764626446
transform -1 0 7807 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_665
timestamp 1764626446
transform -1 0 7807 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_666
timestamp 1764626446
transform -1 0 6499 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_667
timestamp 1764626446
transform -1 0 6499 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_668
timestamp 1764626446
transform -1 0 6499 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_669
timestamp 1764626446
transform -1 0 6499 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_670
timestamp 1764626446
transform -1 0 6499 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_671
timestamp 1764626446
transform -1 0 6499 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_672
timestamp 1764626446
transform -1 0 6499 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_673
timestamp 1764626446
transform -1 0 7807 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_674
timestamp 1764626446
transform -1 0 7371 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_675
timestamp 1764626446
transform -1 0 7371 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_676
timestamp 1764626446
transform -1 0 7371 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_677
timestamp 1764626446
transform -1 0 6063 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_678
timestamp 1764626446
transform -1 0 6063 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_679
timestamp 1764626446
transform -1 0 6063 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_680
timestamp 1764626446
transform -1 0 6063 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_681
timestamp 1764626446
transform -1 0 6063 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_682
timestamp 1764626446
transform -1 0 6063 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_683
timestamp 1764626446
transform -1 0 6063 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_684
timestamp 1764626446
transform -1 0 7371 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_685
timestamp 1764626446
transform -1 0 7371 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_686
timestamp 1764626446
transform -1 0 5627 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_687
timestamp 1764626446
transform -1 0 5627 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_688
timestamp 1764626446
transform 1 0 1119 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_689
timestamp 1764626446
transform 1 0 1119 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_690
timestamp 1764626446
transform 1 0 1555 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_691
timestamp 1764626446
transform 1 0 1555 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_692
timestamp 1764626446
transform -1 0 5191 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_693
timestamp 1764626446
transform -1 0 5191 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_694
timestamp 1764626446
transform -1 0 4755 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_695
timestamp 1764626446
transform -1 0 4755 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_696
timestamp 1764626446
transform -1 0 6935 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_697
timestamp 1764626446
transform -1 0 6935 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_698
timestamp 1764626446
transform -1 0 6499 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_699
timestamp 1764626446
transform -1 0 6499 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_700
timestamp 1764626446
transform 1 0 2863 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_701
timestamp 1764626446
transform 1 0 2863 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_702
timestamp 1764626446
transform -1 0 6063 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_703
timestamp 1764626446
transform -1 0 6063 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_704
timestamp 1764626446
transform -1 0 5627 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_705
timestamp 1764626446
transform -1 0 5627 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_706
timestamp 1764626446
transform -1 0 7807 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_707
timestamp 1764626446
transform -1 0 7807 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_708
timestamp 1764626446
transform -1 0 7371 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_709
timestamp 1764626446
transform -1 0 7371 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_710
timestamp 1764626446
transform 1 0 3299 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_711
timestamp 1764626446
transform 1 0 3299 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_712
timestamp 1764626446
transform 1 0 1991 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_713
timestamp 1764626446
transform 1 0 1991 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_714
timestamp 1764626446
transform 1 0 2427 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_715
timestamp 1764626446
transform 1 0 2427 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_716
timestamp 1764626446
transform 1 0 247 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_717
timestamp 1764626446
transform 1 0 247 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_718
timestamp 1764626446
transform 1 0 683 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_719
timestamp 1764626446
transform 1 0 683 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_720
timestamp 1764626446
transform -1 0 12571 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_721
timestamp 1764626446
transform -1 0 15187 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_722
timestamp 1764626446
transform -1 0 13007 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_723
timestamp 1764626446
transform -1 0 13443 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_724
timestamp 1764626446
transform -1 0 14751 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_725
timestamp 1764626446
transform -1 0 14751 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_726
timestamp 1764626446
transform -1 0 14315 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_727
timestamp 1764626446
transform -1 0 14315 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_728
timestamp 1764626446
transform -1 0 13007 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_729
timestamp 1764626446
transform -1 0 13007 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_730
timestamp 1764626446
transform -1 0 13007 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_731
timestamp 1764626446
transform -1 0 13007 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_732
timestamp 1764626446
transform -1 0 13443 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_733
timestamp 1764626446
transform -1 0 13443 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_734
timestamp 1764626446
transform -1 0 13443 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_735
timestamp 1764626446
transform -1 0 13443 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_736
timestamp 1764626446
transform -1 0 13007 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_737
timestamp 1764626446
transform -1 0 15187 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_738
timestamp 1764626446
transform -1 0 12571 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_739
timestamp 1764626446
transform -1 0 12571 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_740
timestamp 1764626446
transform -1 0 12571 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_741
timestamp 1764626446
transform -1 0 12571 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_742
timestamp 1764626446
transform -1 0 12571 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_743
timestamp 1764626446
transform -1 0 15187 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_744
timestamp 1764626446
transform -1 0 15187 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_745
timestamp 1764626446
transform -1 0 15187 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_746
timestamp 1764626446
transform -1 0 15187 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_747
timestamp 1764626446
transform -1 0 13443 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_748
timestamp 1764626446
transform -1 0 14315 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_749
timestamp 1764626446
transform -1 0 13879 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_750
timestamp 1764626446
transform -1 0 14315 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_751
timestamp 1764626446
transform -1 0 14751 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_752
timestamp 1764626446
transform -1 0 13879 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_753
timestamp 1764626446
transform -1 0 13879 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_754
timestamp 1764626446
transform -1 0 13879 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_755
timestamp 1764626446
transform -1 0 13879 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_756
timestamp 1764626446
transform -1 0 13879 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_757
timestamp 1764626446
transform -1 0 14315 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_758
timestamp 1764626446
transform -1 0 14315 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_759
timestamp 1764626446
transform -1 0 15623 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_760
timestamp 1764626446
transform -1 0 14751 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_761
timestamp 1764626446
transform -1 0 14751 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_762
timestamp 1764626446
transform -1 0 15623 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_763
timestamp 1764626446
transform -1 0 15623 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_764
timestamp 1764626446
transform -1 0 15623 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_765
timestamp 1764626446
transform -1 0 15623 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_766
timestamp 1764626446
transform -1 0 15623 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_767
timestamp 1764626446
transform -1 0 14751 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_768
timestamp 1764626446
transform 1 0 10679 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_769
timestamp 1764626446
transform 1 0 8063 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_770
timestamp 1764626446
transform 1 0 10679 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_771
timestamp 1764626446
transform 1 0 10679 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_772
timestamp 1764626446
transform 1 0 9807 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_773
timestamp 1764626446
transform 1 0 9807 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_774
timestamp 1764626446
transform 1 0 8935 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_775
timestamp 1764626446
transform 1 0 8935 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_776
timestamp 1764626446
transform 1 0 8935 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_777
timestamp 1764626446
transform 1 0 8935 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_778
timestamp 1764626446
transform 1 0 8063 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_779
timestamp 1764626446
transform 1 0 8935 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_780
timestamp 1764626446
transform 1 0 9371 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_781
timestamp 1764626446
transform 1 0 9371 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_782
timestamp 1764626446
transform 1 0 11115 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_783
timestamp 1764626446
transform 1 0 11115 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_784
timestamp 1764626446
transform 1 0 11115 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_785
timestamp 1764626446
transform 1 0 11115 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_786
timestamp 1764626446
transform 1 0 11115 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_787
timestamp 1764626446
transform 1 0 9371 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_788
timestamp 1764626446
transform 1 0 8063 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_789
timestamp 1764626446
transform 1 0 8063 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_790
timestamp 1764626446
transform 1 0 8063 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_791
timestamp 1764626446
transform 1 0 8063 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_792
timestamp 1764626446
transform 1 0 9371 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_793
timestamp 1764626446
transform 1 0 8935 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_794
timestamp 1764626446
transform 1 0 9371 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_795
timestamp 1764626446
transform 1 0 10243 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_796
timestamp 1764626446
transform 1 0 10243 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_797
timestamp 1764626446
transform 1 0 10243 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_798
timestamp 1764626446
transform 1 0 10243 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_799
timestamp 1764626446
transform 1 0 10243 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_800
timestamp 1764626446
transform 1 0 9807 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_801
timestamp 1764626446
transform 1 0 8499 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_802
timestamp 1764626446
transform 1 0 8499 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_803
timestamp 1764626446
transform 1 0 8499 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_804
timestamp 1764626446
transform 1 0 9807 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_805
timestamp 1764626446
transform 1 0 9807 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_806
timestamp 1764626446
transform 1 0 9807 0 1 24240
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_807
timestamp 1764626446
transform 1 0 10243 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_808
timestamp 1764626446
transform 1 0 9371 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_809
timestamp 1764626446
transform 1 0 8499 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_810
timestamp 1764626446
transform 1 0 11115 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_811
timestamp 1764626446
transform 1 0 10679 0 1 20604
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_812
timestamp 1764626446
transform 1 0 10679 0 1 21816
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_813
timestamp 1764626446
transform 1 0 8499 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_814
timestamp 1764626446
transform 1 0 8499 0 1 26664
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_815
timestamp 1764626446
transform 1 0 10679 0 1 23028
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_816
timestamp 1764626446
transform 1 0 8499 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_817
timestamp 1764626446
transform 1 0 8499 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_818
timestamp 1764626446
transform 1 0 8935 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_819
timestamp 1764626446
transform 1 0 10679 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_820
timestamp 1764626446
transform 1 0 10679 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_821
timestamp 1764626446
transform 1 0 10679 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_822
timestamp 1764626446
transform 1 0 10679 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_823
timestamp 1764626446
transform 1 0 10679 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_824
timestamp 1764626446
transform 1 0 10679 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_825
timestamp 1764626446
transform 1 0 10679 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_826
timestamp 1764626446
transform 1 0 8935 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_827
timestamp 1764626446
transform 1 0 8499 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_828
timestamp 1764626446
transform 1 0 8499 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_829
timestamp 1764626446
transform 1 0 8935 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_830
timestamp 1764626446
transform 1 0 11115 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_831
timestamp 1764626446
transform 1 0 11115 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_832
timestamp 1764626446
transform 1 0 11115 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_833
timestamp 1764626446
transform 1 0 11115 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_834
timestamp 1764626446
transform 1 0 11115 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_835
timestamp 1764626446
transform 1 0 11115 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_836
timestamp 1764626446
transform 1 0 8063 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_837
timestamp 1764626446
transform 1 0 8063 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_838
timestamp 1764626446
transform 1 0 8063 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_839
timestamp 1764626446
transform 1 0 8063 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_840
timestamp 1764626446
transform 1 0 8063 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_841
timestamp 1764626446
transform 1 0 8063 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_842
timestamp 1764626446
transform 1 0 8063 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_843
timestamp 1764626446
transform 1 0 11115 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_844
timestamp 1764626446
transform 1 0 8935 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_845
timestamp 1764626446
transform 1 0 8499 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_846
timestamp 1764626446
transform 1 0 8499 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_847
timestamp 1764626446
transform 1 0 8935 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_848
timestamp 1764626446
transform 1 0 9807 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_849
timestamp 1764626446
transform 1 0 9807 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_850
timestamp 1764626446
transform 1 0 9807 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_851
timestamp 1764626446
transform 1 0 9807 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_852
timestamp 1764626446
transform 1 0 9807 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_853
timestamp 1764626446
transform 1 0 9807 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_854
timestamp 1764626446
transform 1 0 9807 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_855
timestamp 1764626446
transform 1 0 9371 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_856
timestamp 1764626446
transform 1 0 8499 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_857
timestamp 1764626446
transform 1 0 9371 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_858
timestamp 1764626446
transform 1 0 9371 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_859
timestamp 1764626446
transform 1 0 9371 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_860
timestamp 1764626446
transform 1 0 10243 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_861
timestamp 1764626446
transform 1 0 10243 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_862
timestamp 1764626446
transform 1 0 10243 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_863
timestamp 1764626446
transform 1 0 10243 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_864
timestamp 1764626446
transform 1 0 10243 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_865
timestamp 1764626446
transform 1 0 10243 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_866
timestamp 1764626446
transform 1 0 10243 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_867
timestamp 1764626446
transform 1 0 9371 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_868
timestamp 1764626446
transform 1 0 9371 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_869
timestamp 1764626446
transform 1 0 9371 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_870
timestamp 1764626446
transform 1 0 8935 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_871
timestamp 1764626446
transform 1 0 8935 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_872
timestamp 1764626446
transform -1 0 13007 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_873
timestamp 1764626446
transform -1 0 13007 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_874
timestamp 1764626446
transform -1 0 13007 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_875
timestamp 1764626446
transform -1 0 13007 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_876
timestamp 1764626446
transform -1 0 13007 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_877
timestamp 1764626446
transform -1 0 13007 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_878
timestamp 1764626446
transform -1 0 13007 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_879
timestamp 1764626446
transform -1 0 14315 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_880
timestamp 1764626446
transform -1 0 14315 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_881
timestamp 1764626446
transform -1 0 14315 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_882
timestamp 1764626446
transform -1 0 14315 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_883
timestamp 1764626446
transform -1 0 12571 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_884
timestamp 1764626446
transform -1 0 12571 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_885
timestamp 1764626446
transform -1 0 12571 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_886
timestamp 1764626446
transform -1 0 12571 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_887
timestamp 1764626446
transform -1 0 12571 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_888
timestamp 1764626446
transform -1 0 12571 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_889
timestamp 1764626446
transform -1 0 12571 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_890
timestamp 1764626446
transform -1 0 14315 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_891
timestamp 1764626446
transform -1 0 15623 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_892
timestamp 1764626446
transform -1 0 15623 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_893
timestamp 1764626446
transform -1 0 15623 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_894
timestamp 1764626446
transform -1 0 15623 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_895
timestamp 1764626446
transform -1 0 15623 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_896
timestamp 1764626446
transform -1 0 15623 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_897
timestamp 1764626446
transform -1 0 15623 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_898
timestamp 1764626446
transform -1 0 15187 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_899
timestamp 1764626446
transform -1 0 15187 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_900
timestamp 1764626446
transform -1 0 15187 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_901
timestamp 1764626446
transform -1 0 15187 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_902
timestamp 1764626446
transform -1 0 15187 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_903
timestamp 1764626446
transform -1 0 15187 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_904
timestamp 1764626446
transform -1 0 15187 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_905
timestamp 1764626446
transform -1 0 13879 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_906
timestamp 1764626446
transform -1 0 13879 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_907
timestamp 1764626446
transform -1 0 13879 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_908
timestamp 1764626446
transform -1 0 13879 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_909
timestamp 1764626446
transform -1 0 13879 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_910
timestamp 1764626446
transform -1 0 13879 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_911
timestamp 1764626446
transform -1 0 13879 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_912
timestamp 1764626446
transform -1 0 13443 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_913
timestamp 1764626446
transform -1 0 13443 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_914
timestamp 1764626446
transform -1 0 13443 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_915
timestamp 1764626446
transform -1 0 13443 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_916
timestamp 1764626446
transform -1 0 13443 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_917
timestamp 1764626446
transform -1 0 13443 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_918
timestamp 1764626446
transform -1 0 13443 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_919
timestamp 1764626446
transform -1 0 14751 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_920
timestamp 1764626446
transform -1 0 14751 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_921
timestamp 1764626446
transform -1 0 14751 0 1 32724
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_922
timestamp 1764626446
transform -1 0 14751 0 1 33936
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_923
timestamp 1764626446
transform -1 0 14751 0 1 35148
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_924
timestamp 1764626446
transform -1 0 14751 0 1 36360
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_925
timestamp 1764626446
transform -1 0 14751 0 1 37572
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_926
timestamp 1764626446
transform -1 0 14315 0 1 30300
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_927
timestamp 1764626446
transform -1 0 14315 0 1 31512
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_928
timestamp 1764626446
transform -1 0 13007 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_929
timestamp 1764626446
transform -1 0 13007 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_930
timestamp 1764626446
transform -1 0 12571 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_931
timestamp 1764626446
transform -1 0 12571 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_932
timestamp 1764626446
transform 1 0 8063 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_933
timestamp 1764626446
transform 1 0 8063 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_934
timestamp 1764626446
transform -1 0 15623 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_935
timestamp 1764626446
transform -1 0 15623 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_936
timestamp 1764626446
transform -1 0 15187 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_937
timestamp 1764626446
transform -1 0 15187 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_938
timestamp 1764626446
transform 1 0 8499 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_939
timestamp 1764626446
transform 1 0 8499 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_940
timestamp 1764626446
transform -1 0 13879 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_941
timestamp 1764626446
transform -1 0 13879 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_942
timestamp 1764626446
transform -1 0 13443 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_943
timestamp 1764626446
transform -1 0 13443 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_944
timestamp 1764626446
transform -1 0 14751 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_945
timestamp 1764626446
transform -1 0 14751 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_946
timestamp 1764626446
transform -1 0 14315 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_947
timestamp 1764626446
transform -1 0 14315 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_948
timestamp 1764626446
transform 1 0 10679 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_949
timestamp 1764626446
transform 1 0 10679 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_950
timestamp 1764626446
transform 1 0 11115 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_951
timestamp 1764626446
transform 1 0 11115 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_952
timestamp 1764626446
transform 1 0 9807 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_953
timestamp 1764626446
transform 1 0 9807 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_954
timestamp 1764626446
transform 1 0 10243 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_955
timestamp 1764626446
transform 1 0 10243 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_956
timestamp 1764626446
transform 1 0 8935 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_957
timestamp 1764626446
transform 1 0 8935 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_958
timestamp 1764626446
transform 1 0 9371 0 1 27876
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_959
timestamp 1764626446
transform 1 0 9371 0 1 29088
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_960
timestamp 1764626446
transform -1 0 13007 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_961
timestamp 1764626446
transform -1 0 13007 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_962
timestamp 1764626446
transform -1 0 12571 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_963
timestamp 1764626446
transform -1 0 12571 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_964
timestamp 1764626446
transform -1 0 5191 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_965
timestamp 1764626446
transform -1 0 5191 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_966
timestamp 1764626446
transform -1 0 4755 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_967
timestamp 1764626446
transform -1 0 4755 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_968
timestamp 1764626446
transform -1 0 6935 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_969
timestamp 1764626446
transform -1 0 6935 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_970
timestamp 1764626446
transform -1 0 6499 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_971
timestamp 1764626446
transform -1 0 6499 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_972
timestamp 1764626446
transform -1 0 6063 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_973
timestamp 1764626446
transform -1 0 6063 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_974
timestamp 1764626446
transform -1 0 5627 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_975
timestamp 1764626446
transform -1 0 5627 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_976
timestamp 1764626446
transform -1 0 7807 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_977
timestamp 1764626446
transform -1 0 7807 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_978
timestamp 1764626446
transform -1 0 7371 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_979
timestamp 1764626446
transform -1 0 7371 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_980
timestamp 1764626446
transform -1 0 15623 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_981
timestamp 1764626446
transform -1 0 15623 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_982
timestamp 1764626446
transform -1 0 15187 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_983
timestamp 1764626446
transform -1 0 15187 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_984
timestamp 1764626446
transform -1 0 13879 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_985
timestamp 1764626446
transform -1 0 13879 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_986
timestamp 1764626446
transform -1 0 13443 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_987
timestamp 1764626446
transform -1 0 13443 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_988
timestamp 1764626446
transform -1 0 14751 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_989
timestamp 1764626446
transform -1 0 14751 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_990
timestamp 1764626446
transform -1 0 14315 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_991
timestamp 1764626446
transform -1 0 14315 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_992
timestamp 1764626446
transform 1 0 1119 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_993
timestamp 1764626446
transform 1 0 1119 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_994
timestamp 1764626446
transform 1 0 1555 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_995
timestamp 1764626446
transform 1 0 1555 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_996
timestamp 1764626446
transform 1 0 2863 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_997
timestamp 1764626446
transform 1 0 2863 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_998
timestamp 1764626446
transform 1 0 3299 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_999
timestamp 1764626446
transform 1 0 3299 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1000
timestamp 1764626446
transform 1 0 1991 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1001
timestamp 1764626446
transform 1 0 1991 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1002
timestamp 1764626446
transform 1 0 2427 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1003
timestamp 1764626446
transform 1 0 2427 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1004
timestamp 1764626446
transform 1 0 247 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1005
timestamp 1764626446
transform 1 0 247 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1006
timestamp 1764626446
transform 1 0 683 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1007
timestamp 1764626446
transform 1 0 683 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1008
timestamp 1764626446
transform 1 0 10679 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1009
timestamp 1764626446
transform 1 0 10679 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1010
timestamp 1764626446
transform 1 0 11115 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1011
timestamp 1764626446
transform 1 0 11115 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1012
timestamp 1764626446
transform 1 0 9807 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1013
timestamp 1764626446
transform 1 0 9807 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1014
timestamp 1764626446
transform 1 0 10243 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1015
timestamp 1764626446
transform 1 0 10243 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1016
timestamp 1764626446
transform 1 0 8935 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1017
timestamp 1764626446
transform 1 0 8935 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1018
timestamp 1764626446
transform 1 0 9371 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1019
timestamp 1764626446
transform 1 0 9371 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1020
timestamp 1764626446
transform 1 0 8063 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1021
timestamp 1764626446
transform 1 0 8063 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1022
timestamp 1764626446
transform 1 0 8499 0 1 18180
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1023
timestamp 1764626446
transform 1 0 8499 0 1 19392
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1024
timestamp 1764626446
transform -1 0 5627 0 1 25452
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1025
timestamp 1764626446
transform -1 0 14751 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1026
timestamp 1764626446
transform -1 0 15187 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1027
timestamp 1764626446
transform -1 0 13879 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1028
timestamp 1764626446
transform -1 0 14315 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1029
timestamp 1764626446
transform -1 0 12571 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1030
timestamp 1764626446
transform -1 0 13007 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1031
timestamp 1764626446
transform -1 0 13443 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1032
timestamp 1764626446
transform 1 0 11115 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1033
timestamp 1764626446
transform 1 0 10243 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1034
timestamp 1764626446
transform 1 0 10679 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1035
timestamp 1764626446
transform 1 0 9371 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1036
timestamp 1764626446
transform 1 0 9807 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1037
timestamp 1764626446
transform 1 0 8499 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1038
timestamp 1764626446
transform 1 0 8935 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1039
timestamp 1764626446
transform 1 0 8063 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1040
timestamp 1764626446
transform -1 0 7371 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1041
timestamp 1764626446
transform -1 0 7807 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1042
timestamp 1764626446
transform -1 0 6499 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1043
timestamp 1764626446
transform -1 0 6935 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1044
timestamp 1764626446
transform -1 0 6063 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1045
timestamp 1764626446
transform -1 0 5627 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1046
timestamp 1764626446
transform -1 0 5191 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1047
timestamp 1764626446
transform -1 0 4755 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1048
timestamp 1764626446
transform 1 0 2863 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1049
timestamp 1764626446
transform 1 0 3299 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1050
timestamp 1764626446
transform 1 0 1991 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1051
timestamp 1764626446
transform 1 0 2427 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1052
timestamp 1764626446
transform 1 0 1119 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1053
timestamp 1764626446
transform 1 0 1555 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1054
timestamp 1764626446
transform 1 0 683 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1055
timestamp 1764626446
transform 1 0 247 0 1 38784
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1056
timestamp 1764626446
transform -1 0 15623 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1057
timestamp 1764626446
transform -1 0 14751 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1058
timestamp 1764626446
transform -1 0 15187 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1059
timestamp 1764626446
transform -1 0 13879 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1060
timestamp 1764626446
transform -1 0 14315 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1061
timestamp 1764626446
transform -1 0 13007 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1062
timestamp 1764626446
transform -1 0 13443 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1063
timestamp 1764626446
transform -1 0 12571 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1064
timestamp 1764626446
transform 1 0 11115 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1065
timestamp 1764626446
transform 1 0 10679 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1066
timestamp 1764626446
transform 1 0 10243 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1067
timestamp 1764626446
transform 1 0 9807 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1068
timestamp 1764626446
transform 1 0 9371 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1069
timestamp 1764626446
transform 1 0 8935 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1070
timestamp 1764626446
transform 1 0 8499 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1071
timestamp 1764626446
transform 1 0 8063 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1072
timestamp 1764626446
transform -1 0 7807 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1073
timestamp 1764626446
transform -1 0 7371 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1074
timestamp 1764626446
transform -1 0 6935 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1075
timestamp 1764626446
transform -1 0 6499 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1076
timestamp 1764626446
transform -1 0 6063 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1077
timestamp 1764626446
transform -1 0 5627 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1078
timestamp 1764626446
transform -1 0 5191 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1079
timestamp 1764626446
transform -1 0 4755 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1080
timestamp 1764626446
transform 1 0 2863 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1081
timestamp 1764626446
transform 1 0 3299 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1082
timestamp 1764626446
transform 1 0 1991 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1083
timestamp 1764626446
transform 1 0 2427 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1084
timestamp 1764626446
transform 1 0 1119 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1085
timestamp 1764626446
transform 1 0 1555 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1086
timestamp 1764626446
transform 1 0 683 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1087
timestamp 1764626446
transform 1 0 247 0 1 39996
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1088
timestamp 1764626446
transform -1 0 15623 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1089
timestamp 1764626446
transform -1 0 14751 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1090
timestamp 1764626446
transform -1 0 15187 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1091
timestamp 1764626446
transform -1 0 13879 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1092
timestamp 1764626446
transform -1 0 14315 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1093
timestamp 1764626446
transform -1 0 13007 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1094
timestamp 1764626446
transform -1 0 13443 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1095
timestamp 1764626446
transform -1 0 12571 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1096
timestamp 1764626446
transform 1 0 11115 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1097
timestamp 1764626446
transform 1 0 10679 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1098
timestamp 1764626446
transform 1 0 10243 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1099
timestamp 1764626446
transform 1 0 9807 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1100
timestamp 1764626446
transform 1 0 9371 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1101
timestamp 1764626446
transform 1 0 8935 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1102
timestamp 1764626446
transform 1 0 8499 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1103
timestamp 1764626446
transform 1 0 8063 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1104
timestamp 1764626446
transform -1 0 7807 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1105
timestamp 1764626446
transform -1 0 7371 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1106
timestamp 1764626446
transform -1 0 6935 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1107
timestamp 1764626446
transform -1 0 6499 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1108
timestamp 1764626446
transform -1 0 6063 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1109
timestamp 1764626446
transform -1 0 5627 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1110
timestamp 1764626446
transform -1 0 5191 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1111
timestamp 1764626446
transform -1 0 4755 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1112
timestamp 1764626446
transform 1 0 2863 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1113
timestamp 1764626446
transform 1 0 3299 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1114
timestamp 1764626446
transform 1 0 1991 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1115
timestamp 1764626446
transform 1 0 2427 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1116
timestamp 1764626446
transform 1 0 1119 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1117
timestamp 1764626446
transform 1 0 1555 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1118
timestamp 1764626446
transform 1 0 683 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1119
timestamp 1764626446
transform 1 0 247 0 1 41208
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1120
timestamp 1764626446
transform -1 0 15623 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1121
timestamp 1764626446
transform -1 0 14751 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1122
timestamp 1764626446
transform -1 0 15187 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1123
timestamp 1764626446
transform -1 0 13879 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1124
timestamp 1764626446
transform -1 0 14315 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1125
timestamp 1764626446
transform -1 0 13007 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1126
timestamp 1764626446
transform -1 0 13443 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1127
timestamp 1764626446
transform -1 0 12571 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1128
timestamp 1764626446
transform 1 0 11115 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1129
timestamp 1764626446
transform 1 0 10679 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1130
timestamp 1764626446
transform 1 0 10243 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1131
timestamp 1764626446
transform 1 0 9807 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1132
timestamp 1764626446
transform 1 0 9371 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1133
timestamp 1764626446
transform 1 0 8935 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1134
timestamp 1764626446
transform 1 0 8499 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1135
timestamp 1764626446
transform 1 0 8063 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1136
timestamp 1764626446
transform -1 0 7807 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1137
timestamp 1764626446
transform -1 0 7371 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1138
timestamp 1764626446
transform -1 0 6935 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1139
timestamp 1764626446
transform -1 0 6499 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1140
timestamp 1764626446
transform -1 0 6063 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1141
timestamp 1764626446
transform -1 0 5627 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1142
timestamp 1764626446
transform -1 0 5191 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1143
timestamp 1764626446
transform -1 0 4755 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1144
timestamp 1764626446
transform 1 0 2863 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1145
timestamp 1764626446
transform 1 0 3299 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1146
timestamp 1764626446
transform 1 0 1991 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1147
timestamp 1764626446
transform 1 0 2427 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1148
timestamp 1764626446
transform 1 0 1119 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1149
timestamp 1764626446
transform 1 0 1555 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1150
timestamp 1764626446
transform 1 0 683 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1151
timestamp 1764626446
transform 1 0 247 0 1 42420
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1152
timestamp 1764626446
transform -1 0 15623 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1153
timestamp 1764626446
transform -1 0 14751 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1154
timestamp 1764626446
transform -1 0 15187 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1155
timestamp 1764626446
transform -1 0 13879 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1156
timestamp 1764626446
transform -1 0 14315 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1157
timestamp 1764626446
transform -1 0 13007 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1158
timestamp 1764626446
transform -1 0 13443 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1159
timestamp 1764626446
transform -1 0 12571 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1160
timestamp 1764626446
transform 1 0 11115 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1161
timestamp 1764626446
transform 1 0 10679 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1162
timestamp 1764626446
transform 1 0 10243 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1163
timestamp 1764626446
transform 1 0 9807 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1164
timestamp 1764626446
transform 1 0 9371 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1165
timestamp 1764626446
transform 1 0 8935 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1166
timestamp 1764626446
transform 1 0 8499 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1167
timestamp 1764626446
transform 1 0 8063 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1168
timestamp 1764626446
transform -1 0 7807 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1169
timestamp 1764626446
transform -1 0 7371 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1170
timestamp 1764626446
transform -1 0 6935 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1171
timestamp 1764626446
transform -1 0 6499 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1172
timestamp 1764626446
transform -1 0 6063 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1173
timestamp 1764626446
transform -1 0 5627 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1174
timestamp 1764626446
transform -1 0 5191 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1175
timestamp 1764626446
transform -1 0 4755 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1176
timestamp 1764626446
transform 1 0 2863 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1177
timestamp 1764626446
transform 1 0 3299 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1178
timestamp 1764626446
transform 1 0 1991 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1179
timestamp 1764626446
transform 1 0 2427 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1180
timestamp 1764626446
transform 1 0 1119 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1181
timestamp 1764626446
transform 1 0 1555 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1182
timestamp 1764626446
transform 1 0 683 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1183
timestamp 1764626446
transform 1 0 247 0 1 43632
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1184
timestamp 1764626446
transform -1 0 15623 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1185
timestamp 1764626446
transform -1 0 14751 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1186
timestamp 1764626446
transform -1 0 15187 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1187
timestamp 1764626446
transform -1 0 13879 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1188
timestamp 1764626446
transform -1 0 14315 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1189
timestamp 1764626446
transform -1 0 13007 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1190
timestamp 1764626446
transform -1 0 13443 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1191
timestamp 1764626446
transform -1 0 12571 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1192
timestamp 1764626446
transform 1 0 11115 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1193
timestamp 1764626446
transform 1 0 10679 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1194
timestamp 1764626446
transform 1 0 10243 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1195
timestamp 1764626446
transform 1 0 9807 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1196
timestamp 1764626446
transform 1 0 9371 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1197
timestamp 1764626446
transform 1 0 8935 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1198
timestamp 1764626446
transform 1 0 8499 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1199
timestamp 1764626446
transform 1 0 8063 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1200
timestamp 1764626446
transform -1 0 7807 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1201
timestamp 1764626446
transform -1 0 7371 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1202
timestamp 1764626446
transform -1 0 6935 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1203
timestamp 1764626446
transform -1 0 6499 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1204
timestamp 1764626446
transform -1 0 6063 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1205
timestamp 1764626446
transform -1 0 5627 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1206
timestamp 1764626446
transform -1 0 5191 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1207
timestamp 1764626446
transform -1 0 4755 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1208
timestamp 1764626446
transform 1 0 2863 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1209
timestamp 1764626446
transform 1 0 3299 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1210
timestamp 1764626446
transform 1 0 1991 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1211
timestamp 1764626446
transform 1 0 2427 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1212
timestamp 1764626446
transform 1 0 1119 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1213
timestamp 1764626446
transform 1 0 1555 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1214
timestamp 1764626446
transform 1 0 683 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1215
timestamp 1764626446
transform 1 0 247 0 1 44844
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1216
timestamp 1764626446
transform -1 0 15623 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1217
timestamp 1764626446
transform -1 0 14751 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1218
timestamp 1764626446
transform -1 0 15187 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1219
timestamp 1764626446
transform -1 0 13879 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1220
timestamp 1764626446
transform -1 0 14315 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1221
timestamp 1764626446
transform -1 0 13007 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1222
timestamp 1764626446
transform -1 0 13443 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1223
timestamp 1764626446
transform -1 0 12571 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1224
timestamp 1764626446
transform 1 0 11115 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1225
timestamp 1764626446
transform 1 0 10679 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1226
timestamp 1764626446
transform 1 0 10243 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1227
timestamp 1764626446
transform 1 0 9807 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1228
timestamp 1764626446
transform 1 0 9371 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1229
timestamp 1764626446
transform 1 0 8935 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1230
timestamp 1764626446
transform 1 0 8499 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1231
timestamp 1764626446
transform 1 0 8063 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1232
timestamp 1764626446
transform -1 0 7807 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1233
timestamp 1764626446
transform -1 0 7371 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1234
timestamp 1764626446
transform -1 0 6935 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1235
timestamp 1764626446
transform -1 0 6499 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1236
timestamp 1764626446
transform -1 0 6063 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1237
timestamp 1764626446
transform -1 0 5627 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1238
timestamp 1764626446
transform -1 0 5191 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1239
timestamp 1764626446
transform -1 0 4755 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1240
timestamp 1764626446
transform 1 0 2863 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1241
timestamp 1764626446
transform 1 0 3299 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1242
timestamp 1764626446
transform 1 0 1991 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1243
timestamp 1764626446
transform 1 0 2427 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1244
timestamp 1764626446
transform 1 0 1119 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1245
timestamp 1764626446
transform 1 0 1555 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1246
timestamp 1764626446
transform 1 0 683 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1247
timestamp 1764626446
transform 1 0 247 0 1 46056
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1248
timestamp 1764626446
transform -1 0 15623 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1249
timestamp 1764626446
transform -1 0 14751 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1250
timestamp 1764626446
transform -1 0 15187 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1251
timestamp 1764626446
transform -1 0 13879 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1252
timestamp 1764626446
transform -1 0 14315 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1253
timestamp 1764626446
transform -1 0 13007 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1254
timestamp 1764626446
transform -1 0 13443 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1255
timestamp 1764626446
transform -1 0 12571 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1256
timestamp 1764626446
transform 1 0 11115 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1257
timestamp 1764626446
transform 1 0 10679 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1258
timestamp 1764626446
transform 1 0 10243 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1259
timestamp 1764626446
transform 1 0 9807 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1260
timestamp 1764626446
transform 1 0 9371 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1261
timestamp 1764626446
transform 1 0 8935 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1262
timestamp 1764626446
transform 1 0 8499 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1263
timestamp 1764626446
transform 1 0 8063 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1264
timestamp 1764626446
transform -1 0 7807 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1265
timestamp 1764626446
transform -1 0 7371 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1266
timestamp 1764626446
transform -1 0 6935 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1267
timestamp 1764626446
transform -1 0 6499 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1268
timestamp 1764626446
transform -1 0 6063 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1269
timestamp 1764626446
transform -1 0 5627 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1270
timestamp 1764626446
transform -1 0 5191 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1271
timestamp 1764626446
transform -1 0 4755 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1272
timestamp 1764626446
transform 1 0 2863 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1273
timestamp 1764626446
transform 1 0 3299 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1274
timestamp 1764626446
transform 1 0 1991 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1275
timestamp 1764626446
transform 1 0 2427 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1276
timestamp 1764626446
transform 1 0 1119 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1277
timestamp 1764626446
transform 1 0 1555 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1278
timestamp 1764626446
transform 1 0 683 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1279
timestamp 1764626446
transform 1 0 247 0 1 47268
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1280
timestamp 1764626446
transform -1 0 15623 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1281
timestamp 1764626446
transform -1 0 14751 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1282
timestamp 1764626446
transform -1 0 15187 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1283
timestamp 1764626446
transform -1 0 13879 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1284
timestamp 1764626446
transform -1 0 14315 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1285
timestamp 1764626446
transform -1 0 13007 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1286
timestamp 1764626446
transform -1 0 13443 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1287
timestamp 1764626446
transform -1 0 12571 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1288
timestamp 1764626446
transform 1 0 11115 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1289
timestamp 1764626446
transform 1 0 10679 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1290
timestamp 1764626446
transform 1 0 10243 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1291
timestamp 1764626446
transform 1 0 9807 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1292
timestamp 1764626446
transform 1 0 9371 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1293
timestamp 1764626446
transform 1 0 8935 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1294
timestamp 1764626446
transform 1 0 8499 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1295
timestamp 1764626446
transform 1 0 8063 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1296
timestamp 1764626446
transform -1 0 7807 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1297
timestamp 1764626446
transform -1 0 7371 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1298
timestamp 1764626446
transform -1 0 6935 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1299
timestamp 1764626446
transform -1 0 6499 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1300
timestamp 1764626446
transform -1 0 6063 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1301
timestamp 1764626446
transform -1 0 5627 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1302
timestamp 1764626446
transform -1 0 5191 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1303
timestamp 1764626446
transform -1 0 4755 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1304
timestamp 1764626446
transform 1 0 2863 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1305
timestamp 1764626446
transform 1 0 3299 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1306
timestamp 1764626446
transform 1 0 1991 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1307
timestamp 1764626446
transform 1 0 2427 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1308
timestamp 1764626446
transform 1 0 1119 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1309
timestamp 1764626446
transform 1 0 1555 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1310
timestamp 1764626446
transform 1 0 683 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1311
timestamp 1764626446
transform 1 0 247 0 1 48480
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1312
timestamp 1764626446
transform -1 0 15623 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1313
timestamp 1764626446
transform -1 0 14751 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1314
timestamp 1764626446
transform -1 0 15187 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1315
timestamp 1764626446
transform -1 0 13879 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1316
timestamp 1764626446
transform -1 0 14315 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1317
timestamp 1764626446
transform -1 0 13007 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1318
timestamp 1764626446
transform -1 0 13443 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1319
timestamp 1764626446
transform -1 0 12571 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1320
timestamp 1764626446
transform 1 0 11115 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1321
timestamp 1764626446
transform 1 0 10679 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1322
timestamp 1764626446
transform 1 0 10243 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1323
timestamp 1764626446
transform 1 0 9807 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1324
timestamp 1764626446
transform 1 0 9371 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1325
timestamp 1764626446
transform 1 0 8935 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1326
timestamp 1764626446
transform 1 0 8499 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1327
timestamp 1764626446
transform 1 0 8063 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1328
timestamp 1764626446
transform -1 0 7807 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1329
timestamp 1764626446
transform -1 0 7371 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1330
timestamp 1764626446
transform -1 0 6935 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1331
timestamp 1764626446
transform -1 0 6499 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1332
timestamp 1764626446
transform -1 0 6063 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1333
timestamp 1764626446
transform -1 0 5627 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1334
timestamp 1764626446
transform -1 0 5191 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1335
timestamp 1764626446
transform -1 0 4755 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1336
timestamp 1764626446
transform 1 0 2863 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1337
timestamp 1764626446
transform 1 0 3299 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1338
timestamp 1764626446
transform 1 0 1991 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1339
timestamp 1764626446
transform 1 0 2427 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1340
timestamp 1764626446
transform 1 0 1119 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1341
timestamp 1764626446
transform 1 0 1555 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1342
timestamp 1764626446
transform 1 0 683 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1343
timestamp 1764626446
transform 1 0 247 0 1 49692
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1344
timestamp 1764626446
transform -1 0 15623 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1345
timestamp 1764626446
transform -1 0 14751 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1346
timestamp 1764626446
transform -1 0 15187 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1347
timestamp 1764626446
transform -1 0 13879 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1348
timestamp 1764626446
transform -1 0 14315 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1349
timestamp 1764626446
transform -1 0 13007 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1350
timestamp 1764626446
transform -1 0 13443 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1351
timestamp 1764626446
transform -1 0 12571 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1352
timestamp 1764626446
transform 1 0 11115 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1353
timestamp 1764626446
transform 1 0 10679 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1354
timestamp 1764626446
transform 1 0 10243 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1355
timestamp 1764626446
transform 1 0 9807 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1356
timestamp 1764626446
transform 1 0 9371 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1357
timestamp 1764626446
transform 1 0 8935 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1358
timestamp 1764626446
transform 1 0 8499 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1359
timestamp 1764626446
transform 1 0 8063 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1360
timestamp 1764626446
transform -1 0 7807 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1361
timestamp 1764626446
transform -1 0 7371 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1362
timestamp 1764626446
transform -1 0 6935 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1363
timestamp 1764626446
transform -1 0 6499 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1364
timestamp 1764626446
transform -1 0 6063 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1365
timestamp 1764626446
transform -1 0 5627 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1366
timestamp 1764626446
transform -1 0 5191 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1367
timestamp 1764626446
transform -1 0 4755 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1368
timestamp 1764626446
transform 1 0 2863 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1369
timestamp 1764626446
transform 1 0 3299 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1370
timestamp 1764626446
transform 1 0 1991 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1371
timestamp 1764626446
transform 1 0 2427 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1372
timestamp 1764626446
transform 1 0 1119 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1373
timestamp 1764626446
transform 1 0 1555 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1374
timestamp 1764626446
transform 1 0 683 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1375
timestamp 1764626446
transform 1 0 247 0 1 50904
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1376
timestamp 1764626446
transform -1 0 15623 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1377
timestamp 1764626446
transform -1 0 14751 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1378
timestamp 1764626446
transform -1 0 15187 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1379
timestamp 1764626446
transform -1 0 13879 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1380
timestamp 1764626446
transform -1 0 14315 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1381
timestamp 1764626446
transform -1 0 13007 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1382
timestamp 1764626446
transform -1 0 13443 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1383
timestamp 1764626446
transform -1 0 12571 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1384
timestamp 1764626446
transform 1 0 11115 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1385
timestamp 1764626446
transform 1 0 10679 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1386
timestamp 1764626446
transform 1 0 10243 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1387
timestamp 1764626446
transform 1 0 9807 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1388
timestamp 1764626446
transform 1 0 9371 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1389
timestamp 1764626446
transform 1 0 8935 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1390
timestamp 1764626446
transform 1 0 8499 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1391
timestamp 1764626446
transform 1 0 8063 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1392
timestamp 1764626446
transform -1 0 7807 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1393
timestamp 1764626446
transform -1 0 7371 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1394
timestamp 1764626446
transform -1 0 6935 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1395
timestamp 1764626446
transform -1 0 6499 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1396
timestamp 1764626446
transform -1 0 6063 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1397
timestamp 1764626446
transform -1 0 5627 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1398
timestamp 1764626446
transform -1 0 5191 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1399
timestamp 1764626446
transform -1 0 4755 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1400
timestamp 1764626446
transform 1 0 2863 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1401
timestamp 1764626446
transform 1 0 3299 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1402
timestamp 1764626446
transform 1 0 1991 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1403
timestamp 1764626446
transform 1 0 2427 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1404
timestamp 1764626446
transform 1 0 1119 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1405
timestamp 1764626446
transform 1 0 1555 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1406
timestamp 1764626446
transform 1 0 683 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1407
timestamp 1764626446
transform 1 0 247 0 1 52116
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1408
timestamp 1764626446
transform -1 0 15623 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1409
timestamp 1764626446
transform -1 0 14751 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1410
timestamp 1764626446
transform -1 0 15187 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1411
timestamp 1764626446
transform -1 0 13879 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1412
timestamp 1764626446
transform -1 0 14315 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1413
timestamp 1764626446
transform -1 0 13007 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1414
timestamp 1764626446
transform -1 0 13443 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1415
timestamp 1764626446
transform -1 0 12571 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1416
timestamp 1764626446
transform 1 0 11115 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1417
timestamp 1764626446
transform 1 0 10679 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1418
timestamp 1764626446
transform 1 0 10243 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1419
timestamp 1764626446
transform 1 0 9807 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1420
timestamp 1764626446
transform 1 0 9371 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1421
timestamp 1764626446
transform 1 0 8935 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1422
timestamp 1764626446
transform 1 0 8499 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1423
timestamp 1764626446
transform 1 0 8063 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1424
timestamp 1764626446
transform -1 0 7807 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1425
timestamp 1764626446
transform -1 0 7371 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1426
timestamp 1764626446
transform -1 0 6935 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1427
timestamp 1764626446
transform -1 0 6499 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1428
timestamp 1764626446
transform -1 0 6063 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1429
timestamp 1764626446
transform -1 0 5627 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1430
timestamp 1764626446
transform -1 0 5191 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1431
timestamp 1764626446
transform -1 0 4755 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1432
timestamp 1764626446
transform 1 0 2863 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1433
timestamp 1764626446
transform 1 0 3299 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1434
timestamp 1764626446
transform 1 0 1991 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1435
timestamp 1764626446
transform 1 0 2427 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1436
timestamp 1764626446
transform 1 0 1119 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1437
timestamp 1764626446
transform 1 0 1555 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1438
timestamp 1764626446
transform 1 0 683 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1439
timestamp 1764626446
transform 1 0 247 0 1 53328
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1440
timestamp 1764626446
transform -1 0 15623 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1441
timestamp 1764626446
transform -1 0 14751 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1442
timestamp 1764626446
transform -1 0 15187 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1443
timestamp 1764626446
transform -1 0 13879 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1444
timestamp 1764626446
transform -1 0 14315 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1445
timestamp 1764626446
transform -1 0 13007 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1446
timestamp 1764626446
transform -1 0 13443 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1447
timestamp 1764626446
transform -1 0 12571 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1448
timestamp 1764626446
transform 1 0 11115 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1449
timestamp 1764626446
transform 1 0 10679 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1450
timestamp 1764626446
transform 1 0 10243 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1451
timestamp 1764626446
transform 1 0 9807 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1452
timestamp 1764626446
transform 1 0 9371 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1453
timestamp 1764626446
transform 1 0 8935 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1454
timestamp 1764626446
transform 1 0 8499 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1455
timestamp 1764626446
transform 1 0 8063 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1456
timestamp 1764626446
transform -1 0 7807 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1457
timestamp 1764626446
transform -1 0 7371 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1458
timestamp 1764626446
transform -1 0 6935 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1459
timestamp 1764626446
transform -1 0 6499 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1460
timestamp 1764626446
transform -1 0 6063 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1461
timestamp 1764626446
transform -1 0 5627 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1462
timestamp 1764626446
transform -1 0 5191 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1463
timestamp 1764626446
transform -1 0 4755 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1464
timestamp 1764626446
transform 1 0 2863 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1465
timestamp 1764626446
transform 1 0 3299 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1466
timestamp 1764626446
transform 1 0 1991 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1467
timestamp 1764626446
transform 1 0 2427 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1468
timestamp 1764626446
transform 1 0 1119 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1469
timestamp 1764626446
transform 1 0 1555 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1470
timestamp 1764626446
transform 1 0 683 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1471
timestamp 1764626446
transform 1 0 247 0 1 54540
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1472
timestamp 1764626446
transform -1 0 15623 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1473
timestamp 1764626446
transform -1 0 14751 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1474
timestamp 1764626446
transform -1 0 15187 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1475
timestamp 1764626446
transform -1 0 13879 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1476
timestamp 1764626446
transform -1 0 14315 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1477
timestamp 1764626446
transform -1 0 13007 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1478
timestamp 1764626446
transform -1 0 13443 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1479
timestamp 1764626446
transform -1 0 12571 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1480
timestamp 1764626446
transform 1 0 11115 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1481
timestamp 1764626446
transform 1 0 10679 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1482
timestamp 1764626446
transform 1 0 10243 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1483
timestamp 1764626446
transform 1 0 9807 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1484
timestamp 1764626446
transform 1 0 9371 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1485
timestamp 1764626446
transform 1 0 8935 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1486
timestamp 1764626446
transform 1 0 8499 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1487
timestamp 1764626446
transform 1 0 8063 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1488
timestamp 1764626446
transform -1 0 7807 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1489
timestamp 1764626446
transform -1 0 7371 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1490
timestamp 1764626446
transform -1 0 6935 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1491
timestamp 1764626446
transform -1 0 6499 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1492
timestamp 1764626446
transform -1 0 6063 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1493
timestamp 1764626446
transform -1 0 5627 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1494
timestamp 1764626446
transform -1 0 5191 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1495
timestamp 1764626446
transform -1 0 4755 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1496
timestamp 1764626446
transform 1 0 2863 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1497
timestamp 1764626446
transform 1 0 3299 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1498
timestamp 1764626446
transform 1 0 1991 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1499
timestamp 1764626446
transform 1 0 2427 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1500
timestamp 1764626446
transform 1 0 1119 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1501
timestamp 1764626446
transform 1 0 1555 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1502
timestamp 1764626446
transform 1 0 683 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1503
timestamp 1764626446
transform 1 0 247 0 1 55752
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1504
timestamp 1764626446
transform -1 0 15623 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1505
timestamp 1764626446
transform -1 0 14751 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1506
timestamp 1764626446
transform -1 0 15187 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1507
timestamp 1764626446
transform -1 0 13879 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1508
timestamp 1764626446
transform -1 0 14315 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1509
timestamp 1764626446
transform -1 0 13007 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1510
timestamp 1764626446
transform -1 0 13443 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1511
timestamp 1764626446
transform -1 0 12571 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1512
timestamp 1764626446
transform 1 0 11115 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1513
timestamp 1764626446
transform 1 0 10679 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1514
timestamp 1764626446
transform 1 0 10243 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1515
timestamp 1764626446
transform 1 0 9807 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1516
timestamp 1764626446
transform 1 0 9371 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1517
timestamp 1764626446
transform 1 0 8935 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1518
timestamp 1764626446
transform 1 0 8499 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1519
timestamp 1764626446
transform 1 0 8063 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1520
timestamp 1764626446
transform -1 0 7807 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1521
timestamp 1764626446
transform -1 0 7371 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1522
timestamp 1764626446
transform -1 0 6935 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1523
timestamp 1764626446
transform -1 0 6499 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1524
timestamp 1764626446
transform -1 0 6063 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1525
timestamp 1764626446
transform -1 0 5627 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1526
timestamp 1764626446
transform -1 0 5191 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1527
timestamp 1764626446
transform -1 0 4755 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1528
timestamp 1764626446
transform 1 0 2863 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1529
timestamp 1764626446
transform 1 0 3299 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1530
timestamp 1764626446
transform 1 0 1991 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1531
timestamp 1764626446
transform 1 0 2427 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1532
timestamp 1764626446
transform 1 0 1119 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1533
timestamp 1764626446
transform 1 0 1555 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1534
timestamp 1764626446
transform 1 0 683 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1535
timestamp 1764626446
transform 1 0 247 0 1 56964
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1536
timestamp 1764626446
transform -1 0 15623 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1537
timestamp 1764626446
transform -1 0 14751 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1538
timestamp 1764626446
transform -1 0 15187 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1539
timestamp 1764626446
transform -1 0 13879 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1540
timestamp 1764626446
transform -1 0 14315 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1541
timestamp 1764626446
transform -1 0 13007 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1542
timestamp 1764626446
transform -1 0 13443 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1543
timestamp 1764626446
transform -1 0 12571 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1544
timestamp 1764626446
transform 1 0 11115 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1545
timestamp 1764626446
transform 1 0 10679 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1546
timestamp 1764626446
transform 1 0 10243 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1547
timestamp 1764626446
transform 1 0 9807 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1548
timestamp 1764626446
transform 1 0 9371 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1549
timestamp 1764626446
transform 1 0 8935 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1550
timestamp 1764626446
transform 1 0 8499 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1551
timestamp 1764626446
transform 1 0 8063 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1552
timestamp 1764626446
transform -1 0 7807 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1553
timestamp 1764626446
transform -1 0 7371 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1554
timestamp 1764626446
transform -1 0 6935 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1555
timestamp 1764626446
transform -1 0 6499 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1556
timestamp 1764626446
transform -1 0 6063 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1557
timestamp 1764626446
transform -1 0 5627 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1558
timestamp 1764626446
transform -1 0 5191 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1559
timestamp 1764626446
transform -1 0 4755 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1560
timestamp 1764626446
transform 1 0 2863 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1561
timestamp 1764626446
transform 1 0 3299 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1562
timestamp 1764626446
transform 1 0 1991 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1563
timestamp 1764626446
transform 1 0 2427 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1564
timestamp 1764626446
transform 1 0 1119 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1565
timestamp 1764626446
transform 1 0 1555 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1566
timestamp 1764626446
transform 1 0 683 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1567
timestamp 1764626446
transform 1 0 247 0 1 58176
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1568
timestamp 1764626446
transform -1 0 15623 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1569
timestamp 1764626446
transform -1 0 14751 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1570
timestamp 1764626446
transform -1 0 15187 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1571
timestamp 1764626446
transform -1 0 13879 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1572
timestamp 1764626446
transform -1 0 14315 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1573
timestamp 1764626446
transform -1 0 13007 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1574
timestamp 1764626446
transform -1 0 13443 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1575
timestamp 1764626446
transform -1 0 12571 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1576
timestamp 1764626446
transform 1 0 11115 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1577
timestamp 1764626446
transform 1 0 10679 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1578
timestamp 1764626446
transform 1 0 10243 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1579
timestamp 1764626446
transform 1 0 9807 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1580
timestamp 1764626446
transform 1 0 9371 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1581
timestamp 1764626446
transform 1 0 8935 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1582
timestamp 1764626446
transform 1 0 8499 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1583
timestamp 1764626446
transform 1 0 8063 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1584
timestamp 1764626446
transform -1 0 7807 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1585
timestamp 1764626446
transform -1 0 7371 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1586
timestamp 1764626446
transform -1 0 6935 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1587
timestamp 1764626446
transform -1 0 6499 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1588
timestamp 1764626446
transform -1 0 6063 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1589
timestamp 1764626446
transform -1 0 5627 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1590
timestamp 1764626446
transform -1 0 5191 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1591
timestamp 1764626446
transform -1 0 4755 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1592
timestamp 1764626446
transform 1 0 2863 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1593
timestamp 1764626446
transform 1 0 3299 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1594
timestamp 1764626446
transform 1 0 1991 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1595
timestamp 1764626446
transform 1 0 2427 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1596
timestamp 1764626446
transform 1 0 1119 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1597
timestamp 1764626446
transform 1 0 1555 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1598
timestamp 1764626446
transform 1 0 683 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1599
timestamp 1764626446
transform 1 0 247 0 1 59388
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1600
timestamp 1764626446
transform -1 0 15623 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1601
timestamp 1764626446
transform -1 0 14751 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1602
timestamp 1764626446
transform -1 0 15187 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1603
timestamp 1764626446
transform -1 0 13879 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1604
timestamp 1764626446
transform -1 0 14315 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1605
timestamp 1764626446
transform -1 0 13007 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1606
timestamp 1764626446
transform -1 0 13443 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1607
timestamp 1764626446
transform -1 0 12571 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1608
timestamp 1764626446
transform 1 0 11115 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1609
timestamp 1764626446
transform 1 0 10679 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1610
timestamp 1764626446
transform 1 0 10243 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1611
timestamp 1764626446
transform 1 0 9807 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1612
timestamp 1764626446
transform 1 0 9371 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1613
timestamp 1764626446
transform 1 0 8935 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1614
timestamp 1764626446
transform 1 0 8499 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1615
timestamp 1764626446
transform 1 0 8063 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1616
timestamp 1764626446
transform -1 0 7807 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1617
timestamp 1764626446
transform -1 0 7371 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1618
timestamp 1764626446
transform -1 0 6935 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1619
timestamp 1764626446
transform -1 0 6499 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1620
timestamp 1764626446
transform -1 0 6063 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1621
timestamp 1764626446
transform -1 0 5627 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1622
timestamp 1764626446
transform -1 0 5191 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1623
timestamp 1764626446
transform -1 0 4755 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1624
timestamp 1764626446
transform 1 0 2863 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1625
timestamp 1764626446
transform 1 0 3299 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1626
timestamp 1764626446
transform 1 0 1991 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1627
timestamp 1764626446
transform 1 0 2427 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1628
timestamp 1764626446
transform 1 0 1119 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1629
timestamp 1764626446
transform 1 0 1555 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1630
timestamp 1764626446
transform 1 0 683 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1631
timestamp 1764626446
transform 1 0 247 0 1 60600
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1632
timestamp 1764626446
transform -1 0 15623 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1633
timestamp 1764626446
transform -1 0 14751 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1634
timestamp 1764626446
transform -1 0 15187 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1635
timestamp 1764626446
transform -1 0 13879 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1636
timestamp 1764626446
transform -1 0 14315 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1637
timestamp 1764626446
transform -1 0 13007 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1638
timestamp 1764626446
transform -1 0 13443 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1639
timestamp 1764626446
transform -1 0 12571 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1640
timestamp 1764626446
transform 1 0 11115 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1641
timestamp 1764626446
transform 1 0 10679 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1642
timestamp 1764626446
transform 1 0 10243 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1643
timestamp 1764626446
transform 1 0 9807 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1644
timestamp 1764626446
transform 1 0 9371 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1645
timestamp 1764626446
transform 1 0 8935 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1646
timestamp 1764626446
transform 1 0 8499 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1647
timestamp 1764626446
transform 1 0 8063 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1648
timestamp 1764626446
transform -1 0 7807 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1649
timestamp 1764626446
transform -1 0 7371 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1650
timestamp 1764626446
transform -1 0 6935 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1651
timestamp 1764626446
transform -1 0 6499 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1652
timestamp 1764626446
transform -1 0 6063 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1653
timestamp 1764626446
transform -1 0 5627 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1654
timestamp 1764626446
transform -1 0 5191 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1655
timestamp 1764626446
transform -1 0 4755 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1656
timestamp 1764626446
transform 1 0 2863 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1657
timestamp 1764626446
transform 1 0 3299 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1658
timestamp 1764626446
transform 1 0 1991 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1659
timestamp 1764626446
transform 1 0 2427 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1660
timestamp 1764626446
transform 1 0 1119 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1661
timestamp 1764626446
transform 1 0 1555 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1662
timestamp 1764626446
transform 1 0 683 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1663
timestamp 1764626446
transform 1 0 247 0 1 61812
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1664
timestamp 1764626446
transform -1 0 15623 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1665
timestamp 1764626446
transform -1 0 14751 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1666
timestamp 1764626446
transform -1 0 15187 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1667
timestamp 1764626446
transform -1 0 13879 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1668
timestamp 1764626446
transform -1 0 14315 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1669
timestamp 1764626446
transform -1 0 13007 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1670
timestamp 1764626446
transform -1 0 13443 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1671
timestamp 1764626446
transform -1 0 12571 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1672
timestamp 1764626446
transform 1 0 11115 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1673
timestamp 1764626446
transform 1 0 10679 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1674
timestamp 1764626446
transform 1 0 10243 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1675
timestamp 1764626446
transform 1 0 9807 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1676
timestamp 1764626446
transform 1 0 9371 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1677
timestamp 1764626446
transform 1 0 8935 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1678
timestamp 1764626446
transform 1 0 8499 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1679
timestamp 1764626446
transform 1 0 8063 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1680
timestamp 1764626446
transform -1 0 7807 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1681
timestamp 1764626446
transform -1 0 7371 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1682
timestamp 1764626446
transform -1 0 6935 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1683
timestamp 1764626446
transform -1 0 6499 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1684
timestamp 1764626446
transform -1 0 6063 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1685
timestamp 1764626446
transform -1 0 5627 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1686
timestamp 1764626446
transform -1 0 5191 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1687
timestamp 1764626446
transform -1 0 4755 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1688
timestamp 1764626446
transform 1 0 2863 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1689
timestamp 1764626446
transform 1 0 3299 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1690
timestamp 1764626446
transform 1 0 1991 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1691
timestamp 1764626446
transform 1 0 2427 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1692
timestamp 1764626446
transform 1 0 1119 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1693
timestamp 1764626446
transform 1 0 1555 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1694
timestamp 1764626446
transform 1 0 683 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1695
timestamp 1764626446
transform 1 0 247 0 1 63024
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1696
timestamp 1764626446
transform -1 0 15623 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1697
timestamp 1764626446
transform -1 0 14751 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1698
timestamp 1764626446
transform -1 0 15187 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1699
timestamp 1764626446
transform -1 0 13879 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1700
timestamp 1764626446
transform -1 0 14315 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1701
timestamp 1764626446
transform -1 0 13007 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1702
timestamp 1764626446
transform -1 0 13443 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1703
timestamp 1764626446
transform -1 0 12571 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1704
timestamp 1764626446
transform 1 0 11115 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1705
timestamp 1764626446
transform 1 0 10679 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1706
timestamp 1764626446
transform 1 0 10243 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1707
timestamp 1764626446
transform 1 0 9807 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1708
timestamp 1764626446
transform 1 0 9371 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1709
timestamp 1764626446
transform 1 0 8935 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1710
timestamp 1764626446
transform 1 0 8499 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1711
timestamp 1764626446
transform 1 0 8063 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1712
timestamp 1764626446
transform -1 0 7807 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1713
timestamp 1764626446
transform -1 0 7371 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1714
timestamp 1764626446
transform -1 0 6935 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1715
timestamp 1764626446
transform -1 0 6499 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1716
timestamp 1764626446
transform -1 0 6063 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1717
timestamp 1764626446
transform -1 0 5627 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1718
timestamp 1764626446
transform -1 0 5191 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1719
timestamp 1764626446
transform -1 0 4755 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1720
timestamp 1764626446
transform 1 0 2863 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1721
timestamp 1764626446
transform 1 0 3299 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1722
timestamp 1764626446
transform 1 0 1991 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1723
timestamp 1764626446
transform 1 0 2427 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1724
timestamp 1764626446
transform 1 0 1119 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1725
timestamp 1764626446
transform 1 0 1555 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1726
timestamp 1764626446
transform 1 0 683 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1727
timestamp 1764626446
transform 1 0 247 0 1 64236
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1728
timestamp 1764626446
transform -1 0 15623 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1729
timestamp 1764626446
transform -1 0 14751 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1730
timestamp 1764626446
transform -1 0 15187 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1731
timestamp 1764626446
transform -1 0 13879 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1732
timestamp 1764626446
transform -1 0 14315 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1733
timestamp 1764626446
transform -1 0 13007 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1734
timestamp 1764626446
transform -1 0 13443 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1735
timestamp 1764626446
transform -1 0 12571 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1736
timestamp 1764626446
transform 1 0 11115 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1737
timestamp 1764626446
transform 1 0 10679 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1738
timestamp 1764626446
transform 1 0 10243 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1739
timestamp 1764626446
transform 1 0 9807 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1740
timestamp 1764626446
transform 1 0 9371 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1741
timestamp 1764626446
transform 1 0 8935 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1742
timestamp 1764626446
transform 1 0 8499 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1743
timestamp 1764626446
transform 1 0 8063 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1744
timestamp 1764626446
transform -1 0 7807 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1745
timestamp 1764626446
transform -1 0 7371 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1746
timestamp 1764626446
transform -1 0 6935 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1747
timestamp 1764626446
transform -1 0 6499 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1748
timestamp 1764626446
transform -1 0 6063 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1749
timestamp 1764626446
transform -1 0 5627 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1750
timestamp 1764626446
transform -1 0 5191 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1751
timestamp 1764626446
transform -1 0 4755 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1752
timestamp 1764626446
transform 1 0 2863 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1753
timestamp 1764626446
transform 1 0 3299 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1754
timestamp 1764626446
transform 1 0 1991 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1755
timestamp 1764626446
transform 1 0 2427 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1756
timestamp 1764626446
transform 1 0 1119 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1757
timestamp 1764626446
transform 1 0 1555 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1758
timestamp 1764626446
transform 1 0 683 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1759
timestamp 1764626446
transform 1 0 247 0 1 65448
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1760
timestamp 1764626446
transform -1 0 15623 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1761
timestamp 1764626446
transform -1 0 14751 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1762
timestamp 1764626446
transform -1 0 15187 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1763
timestamp 1764626446
transform -1 0 13879 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1764
timestamp 1764626446
transform -1 0 14315 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1765
timestamp 1764626446
transform -1 0 13007 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1766
timestamp 1764626446
transform -1 0 13443 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1767
timestamp 1764626446
transform -1 0 12571 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1768
timestamp 1764626446
transform 1 0 11115 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1769
timestamp 1764626446
transform 1 0 10679 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1770
timestamp 1764626446
transform 1 0 10243 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1771
timestamp 1764626446
transform 1 0 9807 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1772
timestamp 1764626446
transform 1 0 9371 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1773
timestamp 1764626446
transform 1 0 8935 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1774
timestamp 1764626446
transform 1 0 8499 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1775
timestamp 1764626446
transform 1 0 8063 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1776
timestamp 1764626446
transform -1 0 7807 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1777
timestamp 1764626446
transform -1 0 7371 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1778
timestamp 1764626446
transform -1 0 6935 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1779
timestamp 1764626446
transform -1 0 6499 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1780
timestamp 1764626446
transform -1 0 6063 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1781
timestamp 1764626446
transform -1 0 5627 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1782
timestamp 1764626446
transform -1 0 5191 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1783
timestamp 1764626446
transform -1 0 4755 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1784
timestamp 1764626446
transform 1 0 2863 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1785
timestamp 1764626446
transform 1 0 3299 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1786
timestamp 1764626446
transform 1 0 1991 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1787
timestamp 1764626446
transform 1 0 2427 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1788
timestamp 1764626446
transform 1 0 1119 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1789
timestamp 1764626446
transform 1 0 1555 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1790
timestamp 1764626446
transform 1 0 683 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1791
timestamp 1764626446
transform 1 0 247 0 1 66660
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1792
timestamp 1764626446
transform -1 0 15623 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1793
timestamp 1764626446
transform -1 0 14751 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1794
timestamp 1764626446
transform -1 0 15187 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1795
timestamp 1764626446
transform -1 0 13879 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1796
timestamp 1764626446
transform -1 0 14315 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1797
timestamp 1764626446
transform -1 0 13007 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1798
timestamp 1764626446
transform -1 0 13443 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1799
timestamp 1764626446
transform -1 0 12571 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1800
timestamp 1764626446
transform 1 0 11115 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1801
timestamp 1764626446
transform 1 0 10679 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1802
timestamp 1764626446
transform 1 0 10243 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1803
timestamp 1764626446
transform 1 0 9807 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1804
timestamp 1764626446
transform 1 0 9371 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1805
timestamp 1764626446
transform 1 0 8935 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1806
timestamp 1764626446
transform 1 0 8499 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1807
timestamp 1764626446
transform 1 0 8063 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1808
timestamp 1764626446
transform -1 0 7807 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1809
timestamp 1764626446
transform -1 0 7371 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1810
timestamp 1764626446
transform -1 0 6935 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1811
timestamp 1764626446
transform -1 0 6499 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1812
timestamp 1764626446
transform -1 0 6063 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1813
timestamp 1764626446
transform -1 0 5627 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1814
timestamp 1764626446
transform -1 0 5191 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1815
timestamp 1764626446
transform -1 0 4755 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1816
timestamp 1764626446
transform 1 0 2863 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1817
timestamp 1764626446
transform 1 0 3299 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1818
timestamp 1764626446
transform 1 0 1991 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1819
timestamp 1764626446
transform 1 0 2427 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1820
timestamp 1764626446
transform 1 0 1119 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1821
timestamp 1764626446
transform 1 0 1555 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1822
timestamp 1764626446
transform 1 0 683 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1823
timestamp 1764626446
transform 1 0 247 0 1 67872
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1824
timestamp 1764626446
transform -1 0 15623 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1825
timestamp 1764626446
transform -1 0 14751 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1826
timestamp 1764626446
transform -1 0 15187 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1827
timestamp 1764626446
transform -1 0 13879 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1828
timestamp 1764626446
transform -1 0 14315 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1829
timestamp 1764626446
transform -1 0 13007 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1830
timestamp 1764626446
transform -1 0 13443 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1831
timestamp 1764626446
transform -1 0 12571 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1832
timestamp 1764626446
transform 1 0 11115 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1833
timestamp 1764626446
transform 1 0 10679 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1834
timestamp 1764626446
transform 1 0 10243 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1835
timestamp 1764626446
transform 1 0 9807 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1836
timestamp 1764626446
transform 1 0 9371 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1837
timestamp 1764626446
transform 1 0 8935 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1838
timestamp 1764626446
transform 1 0 8499 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1839
timestamp 1764626446
transform 1 0 8063 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1840
timestamp 1764626446
transform -1 0 7807 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1841
timestamp 1764626446
transform -1 0 7371 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1842
timestamp 1764626446
transform -1 0 6935 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1843
timestamp 1764626446
transform -1 0 6499 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1844
timestamp 1764626446
transform -1 0 6063 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1845
timestamp 1764626446
transform -1 0 5627 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1846
timestamp 1764626446
transform -1 0 5191 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1847
timestamp 1764626446
transform -1 0 4755 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1848
timestamp 1764626446
transform 1 0 2863 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1849
timestamp 1764626446
transform 1 0 3299 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1850
timestamp 1764626446
transform 1 0 1991 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1851
timestamp 1764626446
transform 1 0 2427 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1852
timestamp 1764626446
transform 1 0 1119 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1853
timestamp 1764626446
transform 1 0 1555 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1854
timestamp 1764626446
transform 1 0 683 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1855
timestamp 1764626446
transform 1 0 247 0 1 69084
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1856
timestamp 1764626446
transform -1 0 15623 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1857
timestamp 1764626446
transform -1 0 14751 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1858
timestamp 1764626446
transform -1 0 15187 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1859
timestamp 1764626446
transform -1 0 13879 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1860
timestamp 1764626446
transform -1 0 14315 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1861
timestamp 1764626446
transform -1 0 13007 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1862
timestamp 1764626446
transform -1 0 13443 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1863
timestamp 1764626446
transform -1 0 12571 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1864
timestamp 1764626446
transform 1 0 11115 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1865
timestamp 1764626446
transform 1 0 10679 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1866
timestamp 1764626446
transform 1 0 10243 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1867
timestamp 1764626446
transform 1 0 9807 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1868
timestamp 1764626446
transform 1 0 9371 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1869
timestamp 1764626446
transform 1 0 8935 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1870
timestamp 1764626446
transform 1 0 8499 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1871
timestamp 1764626446
transform 1 0 8063 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1872
timestamp 1764626446
transform -1 0 7807 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1873
timestamp 1764626446
transform -1 0 7371 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1874
timestamp 1764626446
transform -1 0 6935 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1875
timestamp 1764626446
transform -1 0 6499 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1876
timestamp 1764626446
transform -1 0 6063 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1877
timestamp 1764626446
transform -1 0 5627 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1878
timestamp 1764626446
transform -1 0 5191 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1879
timestamp 1764626446
transform -1 0 4755 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1880
timestamp 1764626446
transform 1 0 2863 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1881
timestamp 1764626446
transform 1 0 3299 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1882
timestamp 1764626446
transform 1 0 1991 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1883
timestamp 1764626446
transform 1 0 2427 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1884
timestamp 1764626446
transform 1 0 1119 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1885
timestamp 1764626446
transform 1 0 1555 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1886
timestamp 1764626446
transform 1 0 683 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1887
timestamp 1764626446
transform 1 0 247 0 1 70296
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1888
timestamp 1764626446
transform -1 0 15623 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1889
timestamp 1764626446
transform -1 0 14751 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1890
timestamp 1764626446
transform -1 0 15187 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1891
timestamp 1764626446
transform -1 0 13879 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1892
timestamp 1764626446
transform -1 0 14315 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1893
timestamp 1764626446
transform -1 0 13007 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1894
timestamp 1764626446
transform -1 0 13443 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1895
timestamp 1764626446
transform -1 0 12571 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1896
timestamp 1764626446
transform 1 0 11115 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1897
timestamp 1764626446
transform 1 0 10679 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1898
timestamp 1764626446
transform 1 0 10243 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1899
timestamp 1764626446
transform 1 0 9807 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1900
timestamp 1764626446
transform 1 0 9371 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1901
timestamp 1764626446
transform 1 0 8935 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1902
timestamp 1764626446
transform 1 0 8499 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1903
timestamp 1764626446
transform 1 0 8063 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1904
timestamp 1764626446
transform -1 0 7807 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1905
timestamp 1764626446
transform -1 0 7371 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1906
timestamp 1764626446
transform -1 0 6935 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1907
timestamp 1764626446
transform -1 0 6499 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1908
timestamp 1764626446
transform -1 0 6063 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1909
timestamp 1764626446
transform -1 0 5627 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1910
timestamp 1764626446
transform -1 0 5191 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1911
timestamp 1764626446
transform -1 0 4755 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1912
timestamp 1764626446
transform 1 0 2863 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1913
timestamp 1764626446
transform 1 0 3299 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1914
timestamp 1764626446
transform 1 0 1991 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1915
timestamp 1764626446
transform 1 0 2427 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1916
timestamp 1764626446
transform 1 0 1119 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1917
timestamp 1764626446
transform 1 0 1555 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1918
timestamp 1764626446
transform 1 0 683 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1919
timestamp 1764626446
transform 1 0 247 0 1 71508
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1920
timestamp 1764626446
transform -1 0 15623 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1921
timestamp 1764626446
transform -1 0 14751 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1922
timestamp 1764626446
transform -1 0 15187 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1923
timestamp 1764626446
transform -1 0 13879 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1924
timestamp 1764626446
transform -1 0 14315 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1925
timestamp 1764626446
transform -1 0 13007 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1926
timestamp 1764626446
transform -1 0 13443 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1927
timestamp 1764626446
transform -1 0 12571 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1928
timestamp 1764626446
transform 1 0 11115 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1929
timestamp 1764626446
transform 1 0 10679 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1930
timestamp 1764626446
transform 1 0 10243 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1931
timestamp 1764626446
transform 1 0 9807 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1932
timestamp 1764626446
transform 1 0 9371 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1933
timestamp 1764626446
transform 1 0 8935 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1934
timestamp 1764626446
transform 1 0 8499 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1935
timestamp 1764626446
transform 1 0 8063 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1936
timestamp 1764626446
transform -1 0 7807 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1937
timestamp 1764626446
transform -1 0 7371 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1938
timestamp 1764626446
transform -1 0 6935 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1939
timestamp 1764626446
transform -1 0 6499 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1940
timestamp 1764626446
transform -1 0 6063 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1941
timestamp 1764626446
transform -1 0 5627 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1942
timestamp 1764626446
transform -1 0 5191 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1943
timestamp 1764626446
transform -1 0 4755 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1944
timestamp 1764626446
transform 1 0 2863 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1945
timestamp 1764626446
transform 1 0 3299 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1946
timestamp 1764626446
transform 1 0 1991 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1947
timestamp 1764626446
transform 1 0 2427 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1948
timestamp 1764626446
transform 1 0 1119 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1949
timestamp 1764626446
transform 1 0 1555 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1950
timestamp 1764626446
transform 1 0 683 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1951
timestamp 1764626446
transform 1 0 247 0 1 72720
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1952
timestamp 1764626446
transform -1 0 15623 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1953
timestamp 1764626446
transform -1 0 14751 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1954
timestamp 1764626446
transform -1 0 15187 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1955
timestamp 1764626446
transform -1 0 13879 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1956
timestamp 1764626446
transform -1 0 14315 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1957
timestamp 1764626446
transform -1 0 13007 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1958
timestamp 1764626446
transform -1 0 13443 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1959
timestamp 1764626446
transform -1 0 12571 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1960
timestamp 1764626446
transform 1 0 11115 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1961
timestamp 1764626446
transform 1 0 10679 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1962
timestamp 1764626446
transform 1 0 10243 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1963
timestamp 1764626446
transform 1 0 9807 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1964
timestamp 1764626446
transform 1 0 9371 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1965
timestamp 1764626446
transform 1 0 8935 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1966
timestamp 1764626446
transform 1 0 8499 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1967
timestamp 1764626446
transform 1 0 8063 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1968
timestamp 1764626446
transform -1 0 7807 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1969
timestamp 1764626446
transform -1 0 7371 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1970
timestamp 1764626446
transform -1 0 6935 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1971
timestamp 1764626446
transform -1 0 6499 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1972
timestamp 1764626446
transform -1 0 6063 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1973
timestamp 1764626446
transform -1 0 5627 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1974
timestamp 1764626446
transform -1 0 5191 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1975
timestamp 1764626446
transform -1 0 4755 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1976
timestamp 1764626446
transform 1 0 2863 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1977
timestamp 1764626446
transform 1 0 3299 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1978
timestamp 1764626446
transform 1 0 1991 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1979
timestamp 1764626446
transform 1 0 2427 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1980
timestamp 1764626446
transform 1 0 1119 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1981
timestamp 1764626446
transform 1 0 1555 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1982
timestamp 1764626446
transform 1 0 683 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1983
timestamp 1764626446
transform 1 0 247 0 1 73932
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1984
timestamp 1764626446
transform -1 0 15623 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1985
timestamp 1764626446
transform -1 0 14751 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1986
timestamp 1764626446
transform -1 0 15187 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1987
timestamp 1764626446
transform -1 0 13879 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1988
timestamp 1764626446
transform -1 0 14315 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1989
timestamp 1764626446
transform -1 0 13007 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1990
timestamp 1764626446
transform -1 0 13443 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1991
timestamp 1764626446
transform -1 0 12571 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1992
timestamp 1764626446
transform 1 0 11115 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1993
timestamp 1764626446
transform 1 0 10679 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1994
timestamp 1764626446
transform 1 0 10243 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1995
timestamp 1764626446
transform 1 0 9807 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1996
timestamp 1764626446
transform 1 0 9371 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1997
timestamp 1764626446
transform 1 0 8935 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1998
timestamp 1764626446
transform 1 0 8499 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1999
timestamp 1764626446
transform 1 0 8063 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2000
timestamp 1764626446
transform -1 0 7807 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2001
timestamp 1764626446
transform -1 0 7371 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2002
timestamp 1764626446
transform -1 0 6935 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2003
timestamp 1764626446
transform -1 0 6499 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2004
timestamp 1764626446
transform -1 0 6063 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2005
timestamp 1764626446
transform -1 0 5627 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2006
timestamp 1764626446
transform -1 0 5191 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2007
timestamp 1764626446
transform -1 0 4755 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2008
timestamp 1764626446
transform 1 0 2863 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2009
timestamp 1764626446
transform 1 0 3299 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2010
timestamp 1764626446
transform 1 0 1991 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2011
timestamp 1764626446
transform 1 0 2427 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2012
timestamp 1764626446
transform 1 0 1119 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2013
timestamp 1764626446
transform 1 0 1555 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2014
timestamp 1764626446
transform 1 0 683 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2015
timestamp 1764626446
transform 1 0 247 0 1 75144
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2016
timestamp 1764626446
transform -1 0 15623 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2017
timestamp 1764626446
transform -1 0 14751 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2018
timestamp 1764626446
transform -1 0 15187 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2019
timestamp 1764626446
transform -1 0 13879 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2020
timestamp 1764626446
transform -1 0 14315 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2021
timestamp 1764626446
transform -1 0 13007 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2022
timestamp 1764626446
transform -1 0 13443 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2023
timestamp 1764626446
transform -1 0 12571 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2024
timestamp 1764626446
transform 1 0 11115 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2025
timestamp 1764626446
transform 1 0 10679 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2026
timestamp 1764626446
transform 1 0 10243 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2027
timestamp 1764626446
transform 1 0 9807 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2028
timestamp 1764626446
transform 1 0 9371 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2029
timestamp 1764626446
transform 1 0 8935 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2030
timestamp 1764626446
transform 1 0 8499 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2031
timestamp 1764626446
transform 1 0 8063 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2032
timestamp 1764626446
transform -1 0 7807 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2033
timestamp 1764626446
transform -1 0 7371 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2034
timestamp 1764626446
transform -1 0 6935 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2035
timestamp 1764626446
transform -1 0 6499 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2036
timestamp 1764626446
transform -1 0 6063 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2037
timestamp 1764626446
transform -1 0 5627 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2038
timestamp 1764626446
transform -1 0 5191 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2039
timestamp 1764626446
transform -1 0 4755 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2040
timestamp 1764626446
transform 1 0 2863 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2041
timestamp 1764626446
transform 1 0 3299 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2042
timestamp 1764626446
transform 1 0 1991 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2043
timestamp 1764626446
transform 1 0 2427 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2044
timestamp 1764626446
transform 1 0 1119 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2045
timestamp 1764626446
transform 1 0 1555 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2046
timestamp 1764626446
transform 1 0 683 0 1 76356
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2047
timestamp 1764626446
transform 1 0 247 0 1 76356
box 30 103 570 1445
use 018SRAM_strap1_2x_3v1024x8m81  018SRAM_strap1_2x_3v1024x8m81_0
array 0 0 -420 0 63 1212
timestamp 1764693440
transform -1 0 8236 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_2x_3v1024x8m81  018SRAM_strap1_2x_3v1024x8m81_1
array 0 0 -420 0 63 1212
timestamp 1764693440
transform -1 0 12144 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_2x_3v1024x8m81  018SRAM_strap1_2x_3v1024x8m81_3
array 0 0 -420 0 63 1212
timestamp 1764693440
transform -1 0 4328 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_0
timestamp 1764625442
transform 1 0 15450 0 1 6708
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_1
timestamp 1764625442
transform 1 0 15450 0 -1 9384
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_2
timestamp 1764625442
transform 1 0 15450 0 -1 8172
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_3
timestamp 1764625442
transform 1 0 15450 0 -1 6960
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_4
timestamp 1764625442
transform 1 0 15450 0 -1 5748
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_5
timestamp 1764625442
transform 1 0 15450 0 -1 4536
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_6
timestamp 1764625442
transform 1 0 15450 0 -1 3324
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_7
timestamp 1764625442
transform 1 0 15450 0 -1 2112
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_8
timestamp 1764625442
transform 1 0 15450 0 -1 900
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_9
timestamp 1764625442
transform 1 0 15450 0 1 648
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_10
timestamp 1764625442
transform 1 0 15450 0 1 1860
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_11
timestamp 1764625442
transform 1 0 15450 0 1 3072
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_12
timestamp 1764625442
transform 1 0 15450 0 1 4284
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_13
timestamp 1764625442
transform 1 0 15450 0 1 7920
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_14
timestamp 1764625442
transform 1 0 15450 0 1 5496
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_15
timestamp 1764625442
transform 1 0 15450 0 1 10344
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_16
timestamp 1764625442
transform 1 0 15450 0 1 11556
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_17
timestamp 1764625442
transform 1 0 15450 0 1 12768
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_18
timestamp 1764625442
transform 1 0 15450 0 1 13980
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_19
timestamp 1764625442
transform 1 0 15450 0 1 15192
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_20
timestamp 1764625442
transform 1 0 15450 0 1 16404
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_21
timestamp 1764625442
transform 1 0 15450 0 1 17616
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_22
timestamp 1764625442
transform 1 0 15450 0 -1 19080
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_23
timestamp 1764625442
transform 1 0 15450 0 -1 17868
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_24
timestamp 1764625442
transform 1 0 15450 0 -1 16656
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_25
timestamp 1764625442
transform 1 0 15450 0 -1 15444
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_26
timestamp 1764625442
transform 1 0 15450 0 -1 14232
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_27
timestamp 1764625442
transform 1 0 15450 0 -1 13020
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_28
timestamp 1764625442
transform 1 0 15450 0 -1 11808
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_29
timestamp 1764625442
transform 1 0 15450 0 1 9132
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_30
timestamp 1764625442
transform 1 0 15450 0 -1 10596
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_31
timestamp 1764625442
transform -1 0 420 0 -1 5748
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_32
timestamp 1764625442
transform -1 0 420 0 -1 4536
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_33
timestamp 1764625442
transform -1 0 420 0 -1 3324
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_34
timestamp 1764625442
transform -1 0 420 0 -1 2112
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_35
timestamp 1764625442
transform -1 0 420 0 -1 900
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_36
timestamp 1764625442
transform -1 0 420 0 1 648
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_37
timestamp 1764625442
transform -1 0 420 0 1 1860
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_38
timestamp 1764625442
transform -1 0 420 0 1 3072
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_39
timestamp 1764625442
transform -1 0 420 0 1 4284
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_40
timestamp 1764625442
transform -1 0 420 0 1 5496
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_41
timestamp 1764625442
transform -1 0 420 0 1 6708
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_42
timestamp 1764625442
transform -1 0 420 0 1 7920
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_43
timestamp 1764625442
transform -1 0 420 0 -1 9384
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_44
timestamp 1764625442
transform -1 0 420 0 -1 8172
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_45
timestamp 1764625442
transform -1 0 420 0 -1 6960
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_46
timestamp 1764625442
transform -1 0 420 0 1 16404
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_47
timestamp 1764625442
transform -1 0 420 0 1 17616
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_48
timestamp 1764625442
transform -1 0 420 0 -1 19080
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_49
timestamp 1764625442
transform -1 0 420 0 -1 17868
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_50
timestamp 1764625442
transform -1 0 420 0 1 10344
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_51
timestamp 1764625442
transform -1 0 420 0 1 11556
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_52
timestamp 1764625442
transform -1 0 420 0 1 12768
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_53
timestamp 1764625442
transform -1 0 420 0 1 13980
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_54
timestamp 1764625442
transform -1 0 420 0 1 15192
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_55
timestamp 1764625442
transform -1 0 420 0 -1 16656
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_56
timestamp 1764625442
transform -1 0 420 0 -1 15444
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_57
timestamp 1764625442
transform -1 0 420 0 -1 14232
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_58
timestamp 1764625442
transform -1 0 420 0 -1 13020
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_59
timestamp 1764625442
transform -1 0 420 0 -1 11808
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_60
timestamp 1764625442
transform -1 0 420 0 1 9132
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_61
timestamp 1764625442
transform -1 0 420 0 -1 10596
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_62
timestamp 1764625442
transform -1 0 420 0 1 21252
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_63
timestamp 1764625442
transform -1 0 420 0 1 22464
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_64
timestamp 1764625442
transform -1 0 420 0 1 23676
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_65
timestamp 1764625442
transform -1 0 420 0 -1 22716
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_66
timestamp 1764625442
transform -1 0 420 0 -1 21504
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_67
timestamp 1764625442
transform -1 0 420 0 1 20040
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_68
timestamp 1764625442
transform -1 0 420 0 -1 28776
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_69
timestamp 1764625442
transform -1 0 420 0 -1 27564
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_70
timestamp 1764625442
transform -1 0 420 0 -1 26352
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_71
timestamp 1764625442
transform -1 0 420 0 1 24888
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_72
timestamp 1764625442
transform -1 0 420 0 1 26100
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_73
timestamp 1764625442
transform -1 0 420 0 1 27312
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_74
timestamp 1764625442
transform -1 0 420 0 -1 25140
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_75
timestamp 1764625442
transform -1 0 420 0 -1 23928
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_76
timestamp 1764625442
transform -1 0 420 0 1 37008
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_77
timestamp 1764625442
transform -1 0 420 0 1 38220
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_78
timestamp 1764625442
transform -1 0 420 0 -1 33624
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_79
timestamp 1764625442
transform -1 0 420 0 -1 32412
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_80
timestamp 1764625442
transform -1 0 420 0 -1 37260
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_81
timestamp 1764625442
transform -1 0 420 0 -1 36048
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_82
timestamp 1764625442
transform -1 0 420 0 -1 31200
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_83
timestamp 1764625442
transform -1 0 420 0 -1 38472
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_84
timestamp 1764625442
transform -1 0 420 0 1 29736
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_85
timestamp 1764625442
transform -1 0 420 0 1 30948
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_86
timestamp 1764625442
transform -1 0 420 0 1 32160
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_87
timestamp 1764625442
transform -1 0 420 0 1 33372
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_88
timestamp 1764625442
transform -1 0 420 0 1 34584
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_89
timestamp 1764625442
transform -1 0 420 0 1 35796
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_90
timestamp 1764625442
transform -1 0 420 0 -1 34836
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_91
timestamp 1764625442
transform -1 0 420 0 1 28524
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_92
timestamp 1764625442
transform -1 0 420 0 -1 29988
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_93
timestamp 1764625442
transform 1 0 15450 0 1 23676
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_94
timestamp 1764625442
transform 1 0 15450 0 -1 27564
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_95
timestamp 1764625442
transform 1 0 15450 0 -1 26352
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_96
timestamp 1764625442
transform 1 0 15450 0 -1 25140
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_97
timestamp 1764625442
transform 1 0 15450 0 1 24888
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_98
timestamp 1764625442
transform 1 0 15450 0 -1 23928
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_99
timestamp 1764625442
transform 1 0 15450 0 -1 28776
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_100
timestamp 1764625442
transform 1 0 15450 0 -1 22716
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_101
timestamp 1764625442
transform 1 0 15450 0 -1 21504
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_102
timestamp 1764625442
transform 1 0 15450 0 1 21252
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_103
timestamp 1764625442
transform 1 0 15450 0 1 22464
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_104
timestamp 1764625442
transform 1 0 15450 0 1 20040
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_105
timestamp 1764625442
transform 1 0 15450 0 1 26100
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_106
timestamp 1764625442
transform 1 0 15450 0 1 27312
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_107
timestamp 1764625442
transform 1 0 15450 0 1 38220
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_108
timestamp 1764625442
transform 1 0 15450 0 1 29736
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_109
timestamp 1764625442
transform 1 0 15450 0 1 30948
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_110
timestamp 1764625442
transform 1 0 15450 0 1 32160
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_111
timestamp 1764625442
transform 1 0 15450 0 1 33372
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_112
timestamp 1764625442
transform 1 0 15450 0 1 34584
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_113
timestamp 1764625442
transform 1 0 15450 0 -1 38472
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_114
timestamp 1764625442
transform 1 0 15450 0 -1 37260
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_115
timestamp 1764625442
transform 1 0 15450 0 -1 36048
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_116
timestamp 1764625442
transform 1 0 15450 0 -1 34836
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_117
timestamp 1764625442
transform 1 0 15450 0 -1 33624
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_118
timestamp 1764625442
transform 1 0 15450 0 -1 32412
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_119
timestamp 1764625442
transform 1 0 15450 0 -1 31200
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_120
timestamp 1764625442
transform 1 0 15450 0 1 37008
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_121
timestamp 1764625442
transform 1 0 15450 0 1 35796
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_122
timestamp 1764625442
transform 1 0 15450 0 1 28524
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_123
timestamp 1764625442
transform 1 0 15450 0 -1 29988
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_124
timestamp 1764625442
transform -1 0 420 0 1 18828
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_125
timestamp 1764625442
transform -1 0 420 0 -1 20292
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_126
timestamp 1764625442
transform 1 0 15450 0 -1 20292
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_127
timestamp 1764625442
transform 1 0 15450 0 1 18828
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_128
timestamp 1764625442
transform 1 0 15450 0 1 39432
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_129
timestamp 1764625442
transform 1 0 15450 0 -1 39684
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_130
timestamp 1764625442
transform -1 0 420 0 -1 39684
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_131
timestamp 1764625442
transform -1 0 420 0 1 39432
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_132
timestamp 1764625442
transform -1 0 420 0 -1 40896
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_133
timestamp 1764625442
transform 1 0 15450 0 -1 40896
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_134
timestamp 1764625442
transform 1 0 15450 0 1 40644
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_135
timestamp 1764625442
transform -1 0 420 0 1 40644
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_136
timestamp 1764625442
transform -1 0 420 0 -1 42108
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_137
timestamp 1764625442
transform 1 0 15450 0 -1 42108
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_138
timestamp 1764625442
transform 1 0 15450 0 1 41856
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_139
timestamp 1764625442
transform -1 0 420 0 1 41856
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_140
timestamp 1764625442
transform -1 0 420 0 -1 43320
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_141
timestamp 1764625442
transform 1 0 15450 0 -1 43320
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_142
timestamp 1764625442
transform 1 0 15450 0 1 43068
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_143
timestamp 1764625442
transform -1 0 420 0 1 43068
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_144
timestamp 1764625442
transform -1 0 420 0 -1 44532
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_145
timestamp 1764625442
transform 1 0 15450 0 -1 44532
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_146
timestamp 1764625442
transform 1 0 15450 0 1 44280
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_147
timestamp 1764625442
transform -1 0 420 0 1 44280
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_148
timestamp 1764625442
transform -1 0 420 0 -1 45744
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_149
timestamp 1764625442
transform 1 0 15450 0 -1 45744
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_150
timestamp 1764625442
transform 1 0 15450 0 1 45492
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_151
timestamp 1764625442
transform -1 0 420 0 1 45492
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_152
timestamp 1764625442
transform -1 0 420 0 -1 46956
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_153
timestamp 1764625442
transform 1 0 15450 0 -1 46956
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_154
timestamp 1764625442
transform 1 0 15450 0 1 46704
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_155
timestamp 1764625442
transform -1 0 420 0 1 46704
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_156
timestamp 1764625442
transform -1 0 420 0 -1 48168
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_157
timestamp 1764625442
transform 1 0 15450 0 -1 48168
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_158
timestamp 1764625442
transform 1 0 15450 0 1 47916
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_159
timestamp 1764625442
transform -1 0 420 0 1 47916
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_160
timestamp 1764625442
transform -1 0 420 0 -1 49380
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_161
timestamp 1764625442
transform 1 0 15450 0 -1 49380
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_162
timestamp 1764625442
transform 1 0 15450 0 1 49128
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_163
timestamp 1764625442
transform -1 0 420 0 1 49128
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_164
timestamp 1764625442
transform -1 0 420 0 -1 50592
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_165
timestamp 1764625442
transform 1 0 15450 0 -1 50592
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_166
timestamp 1764625442
transform 1 0 15450 0 1 50340
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_167
timestamp 1764625442
transform -1 0 420 0 1 50340
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_168
timestamp 1764625442
transform -1 0 420 0 -1 51804
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_169
timestamp 1764625442
transform 1 0 15450 0 -1 51804
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_170
timestamp 1764625442
transform 1 0 15450 0 1 51552
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_171
timestamp 1764625442
transform -1 0 420 0 1 51552
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_172
timestamp 1764625442
transform -1 0 420 0 -1 53016
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_173
timestamp 1764625442
transform 1 0 15450 0 -1 53016
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_174
timestamp 1764625442
transform 1 0 15450 0 1 52764
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_175
timestamp 1764625442
transform -1 0 420 0 1 52764
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_176
timestamp 1764625442
transform -1 0 420 0 -1 54228
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_177
timestamp 1764625442
transform 1 0 15450 0 -1 54228
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_178
timestamp 1764625442
transform 1 0 15450 0 1 53976
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_179
timestamp 1764625442
transform -1 0 420 0 1 53976
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_180
timestamp 1764625442
transform -1 0 420 0 -1 55440
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_181
timestamp 1764625442
transform 1 0 15450 0 -1 55440
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_182
timestamp 1764625442
transform 1 0 15450 0 1 55188
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_183
timestamp 1764625442
transform -1 0 420 0 1 55188
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_184
timestamp 1764625442
transform -1 0 420 0 -1 56652
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_185
timestamp 1764625442
transform 1 0 15450 0 -1 56652
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_186
timestamp 1764625442
transform 1 0 15450 0 1 56400
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_187
timestamp 1764625442
transform -1 0 420 0 1 56400
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_188
timestamp 1764625442
transform -1 0 420 0 -1 57864
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_189
timestamp 1764625442
transform 1 0 15450 0 -1 57864
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_190
timestamp 1764625442
transform 1 0 15450 0 1 57612
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_191
timestamp 1764625442
transform -1 0 420 0 1 57612
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_192
timestamp 1764625442
transform -1 0 420 0 -1 59076
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_193
timestamp 1764625442
transform 1 0 15450 0 -1 59076
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_194
timestamp 1764625442
transform 1 0 15450 0 1 58824
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_195
timestamp 1764625442
transform -1 0 420 0 1 58824
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_196
timestamp 1764625442
transform -1 0 420 0 -1 60288
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_197
timestamp 1764625442
transform 1 0 15450 0 -1 60288
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_198
timestamp 1764625442
transform 1 0 15450 0 1 60036
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_199
timestamp 1764625442
transform -1 0 420 0 1 60036
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_200
timestamp 1764625442
transform -1 0 420 0 -1 61500
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_201
timestamp 1764625442
transform 1 0 15450 0 -1 61500
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_202
timestamp 1764625442
transform 1 0 15450 0 1 61248
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_203
timestamp 1764625442
transform -1 0 420 0 1 61248
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_204
timestamp 1764625442
transform -1 0 420 0 -1 62712
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_205
timestamp 1764625442
transform 1 0 15450 0 -1 62712
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_206
timestamp 1764625442
transform 1 0 15450 0 1 62460
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_207
timestamp 1764625442
transform -1 0 420 0 1 62460
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_208
timestamp 1764625442
transform -1 0 420 0 -1 63924
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_209
timestamp 1764625442
transform 1 0 15450 0 -1 63924
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_210
timestamp 1764625442
transform 1 0 15450 0 1 63672
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_211
timestamp 1764625442
transform -1 0 420 0 1 63672
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_212
timestamp 1764625442
transform -1 0 420 0 -1 65136
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_213
timestamp 1764625442
transform 1 0 15450 0 -1 65136
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_214
timestamp 1764625442
transform 1 0 15450 0 1 64884
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_215
timestamp 1764625442
transform -1 0 420 0 1 64884
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_216
timestamp 1764625442
transform -1 0 420 0 -1 66348
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_217
timestamp 1764625442
transform 1 0 15450 0 -1 66348
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_218
timestamp 1764625442
transform 1 0 15450 0 1 66096
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_219
timestamp 1764625442
transform -1 0 420 0 1 66096
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_220
timestamp 1764625442
transform -1 0 420 0 -1 67560
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_221
timestamp 1764625442
transform 1 0 15450 0 -1 67560
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_222
timestamp 1764625442
transform 1 0 15450 0 1 67308
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_223
timestamp 1764625442
transform -1 0 420 0 1 67308
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_224
timestamp 1764625442
transform -1 0 420 0 -1 68772
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_225
timestamp 1764625442
transform 1 0 15450 0 -1 68772
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_226
timestamp 1764625442
transform 1 0 15450 0 1 68520
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_227
timestamp 1764625442
transform -1 0 420 0 1 68520
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_228
timestamp 1764625442
transform -1 0 420 0 -1 69984
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_229
timestamp 1764625442
transform 1 0 15450 0 -1 69984
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_230
timestamp 1764625442
transform 1 0 15450 0 1 69732
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_231
timestamp 1764625442
transform -1 0 420 0 1 69732
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_232
timestamp 1764625442
transform -1 0 420 0 -1 71196
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_233
timestamp 1764625442
transform 1 0 15450 0 -1 71196
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_234
timestamp 1764625442
transform 1 0 15450 0 1 70944
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_235
timestamp 1764625442
transform -1 0 420 0 1 70944
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_236
timestamp 1764625442
transform -1 0 420 0 -1 72408
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_237
timestamp 1764625442
transform 1 0 15450 0 -1 72408
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_238
timestamp 1764625442
transform 1 0 15450 0 1 72156
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_239
timestamp 1764625442
transform -1 0 420 0 1 72156
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_240
timestamp 1764625442
transform -1 0 420 0 -1 73620
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_241
timestamp 1764625442
transform 1 0 15450 0 -1 73620
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_242
timestamp 1764625442
transform 1 0 15450 0 1 73368
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_243
timestamp 1764625442
transform -1 0 420 0 1 73368
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_244
timestamp 1764625442
transform -1 0 420 0 -1 74832
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_245
timestamp 1764625442
transform 1 0 15450 0 -1 74832
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_246
timestamp 1764625442
transform 1 0 15450 0 1 74580
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_247
timestamp 1764625442
transform -1 0 420 0 1 74580
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_248
timestamp 1764625442
transform -1 0 420 0 -1 76044
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_249
timestamp 1764625442
transform 1 0 15450 0 -1 76044
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_250
timestamp 1764625442
transform 1 0 15450 0 1 75792
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_251
timestamp 1764625442
transform -1 0 420 0 1 75792
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_252
timestamp 1764625442
transform -1 0 420 0 -1 77256
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_253
timestamp 1764625442
transform 1 0 15450 0 -1 77256
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_254
timestamp 1764625442
transform 1 0 15450 0 1 77004
box 91 55 511 797
use 018SRAM_strap1_bndry_3v1024x8m81  018SRAM_strap1_bndry_3v1024x8m81_255
timestamp 1764625442
transform -1 0 420 0 1 77004
box 91 55 511 797
<< end >>
