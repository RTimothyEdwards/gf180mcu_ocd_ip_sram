magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< nwell >>
rect -138 -42 -71 132
rect -68 -41 110 132
rect 111 -41 209 132
rect 211 -41 273 132
rect -68 -42 273 -41
rect -138 -63 273 -42
<< polysilicon >>
rect -41 1178 14 1211
rect 118 1178 174 1211
rect -41 -33 14 0
rect 118 -33 174 0
use pmos_5p043105913020100_512x8m81  pmos_5p043105913020100_512x8m81_0
timestamp 1763765945
transform 1 0 -14 0 1 0
box -202 -86 362 1264
<< end >>
