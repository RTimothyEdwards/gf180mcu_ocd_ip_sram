* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

**************************************
* Revision: 1.0
**************************************


*.SCALE METER

.SUBCKT power_route_04
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_PSUB_I01
** N=2765 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_PSUB_I04
** N=3805 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_PSUB$$47122476
** N=5 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nfet_03v3_I12
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pfet_03v3_I13 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
XM0 2 3 1 4 pfet_03v3 L=2.8e-07 W=3.175e-06 AD=2.9964e-12 AS=2.9964e-12 PD=1.45e-05 PS=1.45e-05 NRD=0.0646109 NRS=0.0646109 m=1 nf=1 $X=0 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pmos_1p2$$46889004 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
X0 1 2 3 4 pfet_03v3_I13 $T=-155 0 0 0 $X=-1195 $Y=-620
.ENDS
***************************************
.SUBCKT nfet_03v3_I02 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
XM0 2 3 1 4 nfet_03v3 L=2.8e-07 W=3.175e-06 AD=2.9964e-12 AS=2.9964e-12 PD=1.45e-05 PS=1.45e-05 NRD=0.0646109 NRS=0.0646109 m=1 nf=1 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT nmos_1p2$$47119404 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
X0 1 2 3 4 nfet_03v3_I02 $T=-155 0 0 0 $X=-835 $Y=-620
.ENDS
***************************************
.SUBCKT ypass_gate vss 3 b d bb db ypass pcb vdd
** N=26 EP=9 IP=25 FDC=5
*.SEEDPROM
X2 bb b pcb vdd pfet_03v3_I13 $T=1240 50985 1 0 $X=200 $Y=43555
X3 bb db 3 vdd pfet_03v3_I13 $T=1250 43050 1 0 $X=210 $Y=35620
X4 b d 3 vdd pmos_1p2$$46889004 $T=1405 15300 1 0 $X=-25 $Y=7790
X5 b d ypass vss nmos_1p2$$47119404 $T=1405 24575 1 0 $X=260 $Y=17090
X6 bb db ypass vss nmos_1p2$$47119404 $T=1405 34595 1 0 $X=260 $Y=27110
.ENDS
***************************************
.SUBCKT mux821 1 2 3 4 5 6 7 8 9 13 14 15 16 17 18 19 20 21 22 23
+ 24 25 26 27 28 29 30 31 32 33 42 43 44 45 46 47 48
** N=86 EP=37 IP=165 FDC=48
*.SEEDPROM
XM0 13 42 1 1 nfet_03v3 L=2.8e-07 W=5.3e-07 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=1510 $Y=2370 $D=2
XM1 16 43 1 1 nfet_03v3 L=2.8e-07 W=5.3e-07 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=3750 $Y=2370 $D=2
XM2 19 44 1 1 nfet_03v3 L=2.8e-07 W=5.3e-07 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=7705 $Y=2370 $D=2
XM3 22 45 1 1 nfet_03v3 L=2.8e-07 W=5.3e-07 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=9945 $Y=2370 $D=2
XM4 25 46 1 1 nfet_03v3 L=2.8e-07 W=5.3e-07 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=13895 $Y=2370 $D=2
XM5 28 47 1 1 nfet_03v3 L=2.8e-07 W=5.3e-07 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=16135 $Y=2370 $D=2
XM6 31 48 1 1 nfet_03v3 L=2.8e-07 W=5.3e-07 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=20090 $Y=2370 $D=2
XM7 2 9 1 1 nfet_03v3 L=2.8e-07 W=5.3e-07 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=22330 $Y=2370 $D=2
X10 5 3 7 8 pfet_03v3_I13 $T=23310 51440 1 0 $X=22270 $Y=44010
X11 5 6 2 8 pfet_03v3_I13 $T=23320 43505 1 0 $X=22280 $Y=36075
X12 3 4 2 8 pmos_1p2$$46889004 $T=23475 15755 1 0 $X=22045 $Y=8245
X13 3 4 9 1 nmos_1p2$$47119404 $T=23475 25030 1 0 $X=22330 $Y=17545
X14 5 6 9 1 nmos_1p2$$47119404 $T=23475 35050 1 0 $X=22330 $Y=27565
X15 1 13 15 4 14 6 42 7 8 ypass_gate $T=3490 455 1 180 $X=-1160 $Y=0
X16 1 16 18 4 17 6 43 7 8 ypass_gate $T=3490 455 0 0 $X=2385 $Y=0
X17 1 19 21 4 20 6 44 7 8 ypass_gate $T=9685 455 1 180 $X=5035 $Y=0
X18 1 22 24 4 23 6 45 7 8 ypass_gate $T=9685 455 0 0 $X=8580 $Y=0
X19 1 25 27 4 26 6 46 7 8 ypass_gate $T=15875 455 1 180 $X=11225 $Y=0
X20 1 28 30 4 29 6 47 7 8 ypass_gate $T=15875 455 0 0 $X=14770 $Y=0
X21 1 31 33 4 32 6 48 7 8 ypass_gate $T=22070 455 1 180 $X=17420 $Y=0
.ENDS
***************************************
.SUBCKT pfet_03v3_I18
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_03v3_I13
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_03v3_I14
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$202587180
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_03v3_I16
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pfet_03v3_I15 1 2 3
** N=3 EP=3 IP=0 FDC=1
XM0 2 3 1 1 pfet_03v3 L=2.8e-07 W=1.595e-06 AD=8.892e-13 AS=1.5048e-12 PD=4.46e-06 PS=8.6e-06 NRD=0.304094 NRS=0.51462 m=1 nf=2 $X=0 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pfet_03v3_I04
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_1p2$$202595372
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$202586156
** N=3 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_1p2$$202596396
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pfet_03v3_I11
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_03v3_I19
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT wen_wm1 vss wep 3 4 5 6 7 8 9 10 11 12 13 men vdd wen GWEN 18 19
** N=43 EP=19 IP=113 FDC=31
XM0 3 wen vss vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=1765 $Y=5060 $D=2
XM1 6 men vss vss nfet_03v3 L=2.8e-07 W=6.35e-07 AD=3.562e-13 AS=6.028e-13 PD=1.89e-06 PS=3.62e-06 NRD=0.189781 NRS=0.321168 m=1 nf=1 $X=1765 $Y=8905 $D=2
XM2 vss GWEN 3 vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=2885 $Y=5060 $D=2
XM3 vss vss 6 vss nfet_03v3 L=2.8e-07 W=6.35e-07 AD=6.028e-13 AS=3.562e-13 PD=3.62e-06 PS=1.89e-06 NRD=0.321168 NRS=0.189781 m=1 nf=1 $X=2885 $Y=8905 $D=2
XM4 4 3 vss vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=5125 $Y=4650 $D=2
XM5 5 6 vss vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=5125 $Y=9315 $D=2
XM6 9 6 4 vss nfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=7660 $Y=8385 $D=2
XM7 7 10 vss vss nfet_03v3 L=2.8e-07 W=6.35e-07 AD=6.028e-13 AS=6.028e-13 PD=3.62e-06 PS=3.62e-06 NRD=0.321168 NRS=0.321168 m=1 nf=1 $X=8920 $Y=4240 $D=2
XM8 11 5 9 vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=9970 $Y=9700 $D=2
XM9 vss 12 11 vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=11090 $Y=9700 $D=2
XM10 vss 9 12 vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=13330 $Y=9700 $D=2
XM11 13 12 vss vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=14450 $Y=9700 $D=2
XM12 wep 7 vss vss nfet_03v3 L=2.8e-07 W=1.12e-06 AD=7.68e-13 AS=7.68e-13 PD=5.12e-06 PS=5.12e-06 NRD=1.2 NRS=1.2 m=1 nf=3 $X=12720 $Y=4810 $D=2
XM13 vss 13 8 vss nfet_03v3 L=2.8e-07 W=6.35e-07 AD=6.028e-13 AS=6.028e-13 PD=3.62e-06 PS=3.62e-06 NRD=0.321168 NRS=0.321168 m=1 nf=1 $X=17810 $Y=9290 $D=2
XM14 men 8 10 vss nfet_03v3 L=2.8e-07 W=2.115e-06 AD=1.1804e-12 AS=1.589e-12 PD=5.58e-06 PS=8.21e-06 NRD=0.229075 NRS=0.30837 m=1 nf=2 $X=20050 $Y=8385 $D=2
XM15 vss 13 10 vss nfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=22290 $Y=8385 $D=2
XM16 18 wen vdd vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=1765 $Y=600 $D=8
XM17 19 men vdd vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=1765 $Y=12055 $D=8
XM18 3 GWEN 18 vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=2885 $Y=600 $D=8
XM19 6 vss 19 vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=2885 $Y=12055 $D=8
XM20 4 3 vdd vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=5125 $Y=600 $D=8
XM21 5 6 vdd vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=5125 $Y=12055 $D=8
XM22 9 5 4 vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=1.17084e-12 AS=9.988e-13 PD=4.78598e-06 PS=5.42e-06 NRD=0.22722 NRS=0.193833 m=1 nf=1 $X=7660 $Y=12055 $D=8
XM23 11 6 9 vdd pfet_03v3 L=2.8e-07 W=4.45e-07 AD=-6.87097e-13 AS=-6.48697e-13 PD=-2.78573e-06 PS=-2.70573e-06 NRD=-0.745548 NRS=-0.703882 m=1 nf=1 $X=9395 $Y=12055 $D=8
XM24 vdd 12 11 vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=1.14386e-12 PD=5.42e-06 PS=4.72975e-06 NRD=0.193833 NRS=0.221983 m=1 nf=1 $X=11090 $Y=12055 $D=8
XM25 vdd 9 12 vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=13330 $Y=12055 $D=8
XM26 13 12 vdd vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=14450 $Y=12055 $D=8
XM27 wep 7 vdd vdd pfet_03v3 L=2.8e-07 W=2.8e-06 AD=1.92e-12 AS=1.92e-12 PD=9.92e-06 PS=9.92e-06 NRD=0.48 NRS=0.48 m=1 nf=3 $X=12720 $Y=870 $D=8
XM28 men 13 10 vdd pfet_03v3 L=2.8e-07 W=2.115e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=20050 $Y=12055 $D=8
X48 vdd 7 10 pfet_03v3_I15 $T=8920 2870 1 0 $X=7880 $Y=540
X49 vdd 8 13 pfet_03v3_I15 $T=16690 12625 0 0 $X=15650 $Y=12005
.ENDS
***************************************
.SUBCKT M1_PSUB$$44997676
** N=7 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pfet_03v3_I02
** N=6 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$46286892
** N=5 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_03v3_I10 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
XM0 2 3 1 4 nfet_03v3 L=2.8e-07 W=5.295e-06 AD=3.3596e-12 AS=3.3596e-12 PD=1.658e-05 PS=1.658e-05 NRD=0.651982 NRS=0.651982 m=1 nf=5 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pfet_03v3_I16 1 2 3 4 5
** N=6 EP=5 IP=0 FDC=2
XM0 2 4 1 2 pfet_03v3 L=2.8e-07 W=5.6e-07 AD=3.12e-13 AS=5.28e-13 PD=1.72e-06 PS=3.28e-06 NRD=0.216667 NRS=0.366667 m=1 nf=1 $X=0 $Y=0 $D=8
XM1 3 5 2 2 pfet_03v3 L=2.8e-07 W=5.6e-07 AD=5.28e-13 AS=3.12e-13 PD=3.28e-06 PS=1.72e-06 NRD=0.366667 NRS=0.216667 m=1 nf=1 $X=1120 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nfet_03v3_I17 1 2 3 4 5
** N=5 EP=5 IP=0 FDC=2
XM0 2 4 1 2 nfet_03v3 L=2.8e-07 W=2.8e-07 AD=1.56e-13 AS=2.64e-13 PD=1.12e-06 PS=2.08e-06 NRD=0.433333 NRS=0.733333 m=1 nf=1 $X=0 $Y=0 $D=2
XM1 3 5 2 2 nfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.64e-13 AS=1.56e-13 PD=2.08e-06 PS=1.12e-06 NRD=0.733333 NRS=0.433333 m=1 nf=1 $X=1120 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pmos_1p2$$46285868
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$46281772
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pfet_03v3_I09
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_03v3_I08 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
XM0 2 3 1 4 nfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.64e-13 AS=2.64e-13 PD=2.08e-06 PS=2.08e-06 NRD=0.733333 NRS=0.733333 m=1 nf=1 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT nfet_03v3_I09
** N=6 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sacntl_2 vss 2 pcb 4 5 6 7 8 9 10 11 18 19 20 21 22 23 24 25 26
+ se vdd men
** N=54 EP=23 IP=83 FDC=39
XM0 2 11 vss vss nfet_03v3 L=2.8e-07 W=1.06e-06 AD=5.928e-13 AS=1.0032e-12 PD=3.32e-06 PS=6.32e-06 NRD=0.45614 NRS=0.77193 m=1 nf=2 $X=795 $Y=26115 $D=2
XM1 4 men vss vss nfet_03v3 L=2.8e-07 W=2.66e-06 AD=1.6872e-12 AS=1.6872e-12 PD=9.8e-06 PS=9.8e-06 NRD=1.29825 NRS=1.29825 m=1 nf=5 $X=855 $Y=4275 $D=2
XM2 vss 10 pcb vss nfet_03v3 L=2.8e-07 W=7.415e-06 AD=4.54e-12 AS=4.54e-12 PD=2.216e-05 PS=2.216e-05 NRD=0.881057 NRS=0.881057 m=1 nf=7 $X=1950 $Y=9235 $D=2
XM3 5 4 vss vss nfet_03v3 L=2.8e-07 W=1.33e-06 AD=7.436e-13 AS=1.2584e-12 PD=3.38e-06 PS=6.6e-06 NRD=0.0909091 NRS=0.153846 m=1 nf=1 $X=10910 $Y=8645 $D=2
XM4 6 11 5 vss nfet_03v3 L=2.8e-07 W=1.33e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=12030 $Y=8645 $D=2
XM5 7 19 6 vss nfet_03v3 L=2.8e-07 W=1.33e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=13150 $Y=8645 $D=2
XM6 8 19 7 vss nfet_03v3 L=2.8e-07 W=1.33e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=14270 $Y=8645 $D=2
XM7 9 11 8 vss nfet_03v3 L=2.8e-07 W=1.33e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=15390 $Y=8645 $D=2
XM8 vss 4 9 vss nfet_03v3 L=2.8e-07 W=1.33e-06 AD=1.2584e-12 AS=7.436e-13 PD=6.6e-06 PS=3.38e-06 NRD=0.153846 NRS=0.0909091 m=1 nf=1 $X=16510 $Y=8645 $D=2
XM9 10 7 vss vss nfet_03v3 L=2.8e-07 W=2.435e-06 AD=1.3572e-12 AS=2.2968e-12 PD=6.26e-06 PS=1.22e-05 NRD=0.199234 NRS=0.337165 m=1 nf=2 $X=18750 $Y=8895 $D=2
XM10 11 20 vss vss nfet_03v3 L=2.8e-07 W=6.7e-07 AD=6.336e-13 AS=6.336e-13 PD=3.76e-06 PS=3.76e-06 NRD=0.305556 NRS=0.305556 m=1 nf=1 $X=21255 $Y=4090 $D=2
XM11 se 19 vss vss nfet_03v3 L=2.8e-07 W=4.235e-06 AD=2.3608e-12 AS=3.178e-12 PD=1.116e-05 PS=1.642e-05 NRD=0.45815 NRS=0.61674 m=1 nf=4 $X=19460 $Y=25030 $D=2
XM12 2 11 vdd vdd pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=3.0008e-12 PD=7.86e-06 PS=1.54e-05 NRD=0.152493 NRS=0.258065 m=1 nf=2 $X=795 $Y=20945 $D=8
XM13 4 men vdd vdd pfet_03v3 L=2.8e-07 W=5.295e-06 AD=3.3596e-12 AS=3.3596e-12 PD=1.658e-05 PS=1.658e-05 NRD=0.651982 NRS=0.651982 m=1 nf=5 $X=855 $Y=590 $D=8
XM14 19 2 vdd vdd pfet_03v3 L=2.8e-07 W=3.175e-06 AD=1.7706e-12 AS=2.1792e-12 PD=8.37e-06 PS=1.1e-05 NRD=0.343612 NRS=0.422907 m=1 nf=3 $X=5370 $Y=20990 $D=8
XM15 vdd 4 19 vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=8730 $Y=20990 $D=8
XM16 pcb 10 vdd vdd pfet_03v3 L=2.8e-07 W=1.909e-05 AD=1.0634e-11 AS=1.21023e-11 PD=4.61e-05 PS=4.6818e-05 NRD=0.635697 NRS=0.723472 m=1 nf=10 $X=830 $Y=14055 $D=8
XM17 7 19 vdd vdd pfet_03v3 L=2.8e-07 W=2.115e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.06e-06 PS=9.96e-06 NRD=0.0572687 NRS=0.0969163 m=1 nf=1 $X=14270 $Y=13710 $D=8
XM18 vdd 11 7 vdd pfet_03v3 L=2.8e-07 W=2.115e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=15390 $Y=13710 $D=8
XM19 7 4 vdd vdd pfet_03v3 L=2.8e-07 W=2.115e-06 AD=1.9976e-12 AS=1.1804e-12 PD=9.96e-06 PS=5.06e-06 NRD=0.0969163 NRS=0.0572687 m=1 nf=1 $X=16510 $Y=13710 $D=8
XM20 vdd 25 26 vdd pfet_03v3 L=2.8e-07 W=5.6e-07 AD=5.28e-13 AS=5.28e-13 PD=3.28e-06 PS=3.28e-06 NRD=0.366667 NRS=0.366667 m=1 nf=1 $X=18950 $Y=1670 $D=8
XM21 10 7 vdd vdd pfet_03v3 L=2.8e-07 W=6.355e-06 AD=4.3584e-12 AS=4.3584e-12 PD=2.008e-05 PS=2.008e-05 NRD=0.211454 NRS=0.211454 m=1 nf=3 $X=18750 $Y=13710 $D=8
XM22 se 19 vdd vdd pfet_03v3 L=2.8e-07 W=1.269e-05 AD=7.072e-12 AS=8.0512e-12 PD=3.24e-05 PS=3.856e-05 NRD=0.955882 NRS=1.08824 m=1 nf=10 $X=12740 $Y=20450 $D=8
X23 vdd 11 20 pfet_03v3_I15 $T=21255 985 0 0 $X=20215 $Y=365
X27 vss 18 2 vss nfet_03v3_I10 $T=5370 25030 0 0 $X=4690 $Y=24410
X28 19 18 4 vss nfet_03v3_I10 $T=12415 25030 0 0 $X=11735 $Y=24410
X29 20 vdd 21 4 vss pfet_03v3_I16 $T=8080 1480 0 0 $X=7040 $Y=860
X30 22 vdd 23 21 22 pfet_03v3_I16 $T=11705 1480 0 0 $X=10665 $Y=860
X31 24 vdd 25 23 24 pfet_03v3_I16 $T=15325 1480 0 0 $X=14285 $Y=860
X32 20 vss 21 4 vss nfet_03v3_I17 $T=8080 4420 0 0 $X=7400 $Y=3800
X33 22 vss 23 21 22 nfet_03v3_I17 $T=11705 4420 0 0 $X=11025 $Y=3800
X34 24 vss 25 23 24 nfet_03v3_I17 $T=15325 4420 0 0 $X=14645 $Y=3800
X39 26 vss 25 vss nfet_03v3_I08 $T=18950 4420 0 0 $X=18270 $Y=3800
.ENDS
***************************************
.SUBCKT nfet_03v3_I05
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pfet_03v3_I10
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pfet_03v3_I03
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_03v3_I01
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT outbuf_oe q vss 3 4 5 15 16 17 18 vdd GWE se qp qn 24
** N=66 EP=15 IP=48 FDC=18
XM0 vss 5 q vss nfet_03v3 L=2.8e-07 W=5.935e-06 AD=3.3072e-12 AS=4.0704e-12 PD=1.584e-05 PS=2.08e-05 NRD=0.735849 NRS=0.90566 m=1 nf=6 $X=395 $Y=2665 $D=2
XM1 3 GWE vss vss nfet_03v3 L=2.8e-07 W=7.45e-07 AD=7.04e-13 AS=7.04e-13 PD=4.08e-06 PS=4.08e-06 NRD=0.275 NRS=0.275 m=1 nf=1 $X=8145 $Y=2720 $D=2
XM2 17 3 vss vss nfet_03v3 L=2.8e-07 W=1.025e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=10105 $Y=2700 $D=2
XM3 vss 16 4 vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=13175 $Y=12845 $D=2
XM4 5 15 4 vss nfet_03v3 L=2.8e-07 W=3.175e-06 AD=2.1792e-12 AS=2.1792e-12 PD=1.1e-05 PS=1.1e-05 NRD=0.422907 NRS=0.422907 m=1 nf=3 $X=12455 $Y=2720 $D=2
XM5 vss se 15 vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=17045 $Y=4035 $D=2
XM6 5 qn 18 vss nfet_03v3 L=2.8e-07 W=2.65e-06 AD=1.4768e-12 AS=1.988e-12 PD=6.72e-06 PS=9.92e-06 NRD=0.183099 NRS=0.246479 m=1 nf=2 $X=19905 $Y=1945 $D=2
XM7 vss 3 18 vss nfet_03v3 L=2.8e-07 W=2.65e-06 AD=1.4768e-12 AS=1.988e-12 PD=6.72e-06 PS=9.92e-06 NRD=0.183099 NRS=0.246479 m=1 nf=2 $X=22145 $Y=1945 $D=2
XM8 vdd 5 q vdd pfet_03v3 L=2.8e-07 W=1.058e-05 AD=5.8968e-12 AS=7.2576e-12 PD=2.58e-05 PS=3.408e-05 NRD=0.412698 NRS=0.507937 m=1 nf=6 $X=395 $Y=6190 $D=8
XM9 3 GWE vdd vdd pfet_03v3 L=2.8e-07 W=1.865e-06 AD=1.76e-12 AS=1.76e-12 PD=8.88e-06 PS=8.88e-06 NRD=0.11 NRS=0.11 m=1 nf=1 $X=8145 $Y=6395 $D=8
XM10 17 3 vdd vdd pfet_03v3 L=2.8e-07 W=2.1e-06 AD=1.98e-12 AS=1.98e-12 PD=9.88e-06 PS=9.88e-06 NRD=0.0977778 NRS=0.0977778 m=1 nf=1 $X=10105 $Y=6175 $D=8
XM11 4 16 vdd vdd pfet_03v3 L=2.8e-07 W=1.06e-06 AD=5.928e-13 AS=1.24202e-12 PD=3.32e-06 PS=5.60564e-06 NRD=0.45614 NRS=0.955691 m=1 nf=2 $X=12055 $Y=10310 $D=8
XM12 5 se 4 vdd pfet_03v3 L=2.8e-07 W=3.175e-06 AD=2.1792e-12 AS=2.1792e-12 PD=1.1e-05 PS=1.1e-05 NRD=0.422907 NRS=0.422907 m=1 nf=3 $X=12455 $Y=6395 $D=8
XM13 16 5 vdd vdd pfet_03v3 L=2.8e-07 W=5.6e-07 AD=5.28e-13 AS=7.79385e-13 PD=3.28e-06 PS=2.57436e-06 NRD=0.366667 NRS=0.541239 m=1 nf=1 $X=15085 $Y=10250 $D=8
XM14 vdd se 15 vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=17045 $Y=7030 $D=8
XM15 5 qp 24 vdd pfet_03v3 L=2.8e-07 W=5.29e-06 AD=2.9484e-12 AS=3.969e-12 PD=1.238e-05 PS=1.841e-05 NRD=0.0917108 NRS=0.123457 m=1 nf=2 $X=19680 $Y=6685 $D=8
XM16 vdd 17 24 vdd pfet_03v3 L=2.8e-07 W=5.29e-06 AD=2.9484e-12 AS=3.969e-12 PD=1.238e-05 PS=1.841e-05 NRD=0.0917108 NRS=0.123457 m=1 nf=2 $X=21920 $Y=6685 $D=8
X22 vss 16 5 vss nfet_03v3_I08 $T=15150 13365 1 0 $X=14470 $Y=12145
.ENDS
***************************************
.SUBCKT pmos_1p2$$46887980 1 2 3
** N=3 EP=3 IP=0 FDC=1
XM0 2 3 1 1 pfet_03v3 L=2.8e-07 W=6.35e-06 AD=5.9884e-12 AS=5.9884e-12 PD=2.81e-05 PS=2.81e-05 NRD=0.0323292 NRS=0.0323292 m=1 nf=1 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pmos_1p2$$46273580 1 2 3
** N=3 EP=3 IP=3 FDC=1
XM0 2 3 1 1 pfet_03v3 L=2.8e-07 W=1.06e-06 AD=5.928e-13 AS=1.0032e-12 PD=3.32e-06 PS=6.32e-06 NRD=0.45614 NRS=0.77193 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nmos_1p2$$46883884 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
XM0 2 3 1 4 nfet_03v3 L=2.8e-07 W=5.29e-06 AD=4.9896e-12 AS=4.9896e-12 PD=2.356e-05 PS=2.356e-05 NRD=0.0388007 NRS=0.0388007 m=1 nf=1 $X=-155 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pfet_03v3_I06 1 2 3 4 5 6
** N=6 EP=6 IP=0 FDC=2
XM0 2 4 1 6 pfet_03v3 L=2.8e-07 W=4.45e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=0 $Y=0 $D=8
XM1 3 5 2 6 pfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=1120 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nfet_03v3_I07 1 2 3 4 5 6
** N=6 EP=6 IP=0 FDC=2
XM0 2 4 1 6 nfet_03v3 L=2.8e-07 W=4.45e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=0 $Y=0 $D=2
XM1 3 5 2 6 nfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=1120 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT nmos_1p2$$46563372 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
XM0 2 3 1 4 nfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=-155 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT M1_NWELL_I01
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT din vss 2 3 4 d db 7 8 9 10 11 12 vdd datain men wep
** N=69 EP=16 IP=73 FDC=24
XM0 2 4 vss vss nfet_03v3 L=2.8e-07 W=6.35e-06 AD=5.9884e-12 AS=5.9884e-12 PD=2.81e-05 PS=2.81e-05 NRD=0.0323292 NRS=0.0323292 m=1 nf=1 $X=260 $Y=10430 $D=2
XM1 3 wep vss vss nfet_03v3 L=2.8e-07 W=5.3e-07 AD=7.866e-13 AS=7.923e-13 PD=3.66e-06 PS=3.67e-06 NRD=0.605263 NRS=0.609649 m=1 nf=1 $X=3600 $Y=38320 $D=2
XM2 vss 10 4 vss nfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=11165 $Y=8655 $D=2
XM3 3 wep vdd vdd pfet_03v3 L=2.8e-07 W=1.385e-06 AD=1.13602e-12 AS=1.7523e-12 PD=4.5e-06 PS=8.3e-06 NRD=0.515152 NRS=0.794613 m=1 nf=2 $X=3025 $Y=35440 $D=8
XM4 vdd 2 7 vdd pfet_03v3 L=2.8e-07 W=5.29e-06 AD=4.9896e-12 AS=4.9896e-12 PD=2.356e-05 PS=2.356e-05 NRD=0.0388007 NRS=0.0388007 m=1 nf=1 $X=6980 $Y=26220 $D=8
X5 4 vdd 10 vdd pfet_03v3_I13 $T=11165 455 0 0 $X=10125 $Y=-165
X6 d 2 3 vdd pmos_1p2$$46889004 $T=2655 26220 0 0 $X=1225 $Y=25510
X7 db 7 3 vdd pmos_1p2$$46889004 $T=4895 26220 0 0 $X=3465 $Y=25510
X9 vdd 2 4 pmos_1p2$$46887980 $T=415 26220 0 0 $X=-1015 $Y=25510
X10 vdd 12 men pmos_1p2$$46273580 $T=2920 7175 1 0 $X=1490 $Y=5355
X11 vdd 11 4 pmos_1p2$$46273580 $T=7060 8140 1 0 $X=5630 $Y=6320
X12 d 2 wep vss nmos_1p2$$46883884 $T=2655 12695 0 0 $X=1510 $Y=12010
X13 db 7 wep vss nmos_1p2$$46883884 $T=4895 12695 0 0 $X=3750 $Y=12010
X14 7 vss 2 vss nmos_1p2$$46883884 $T=7135 12695 0 0 $X=5990 $Y=12010
X15 8 vdd 9 datain 8 vdd pfet_03v3_I06 $T=2765 3195 0 0 $X=1725 $Y=2575
X16 9 10 11 men 12 vdd pfet_03v3_I06 $T=6905 3605 0 0 $X=5865 $Y=2985
X17 8 vss 9 datain 8 vss nfet_03v3_I07 $T=2765 1790 1 0 $X=2085 $Y=210
X18 9 10 11 12 men vss nfet_03v3_I07 $T=6905 725 0 0 $X=6225 $Y=105
X19 vss 12 men vss nmos_1p2$$46563372 $T=3470 9035 0 0 $X=2325 $Y=8350
X20 vss 11 4 vss nmos_1p2$$46563372 $T=7060 10495 1 0 $X=5915 $Y=8860
.ENDS
***************************************
.SUBCKT nmos_1p2$$46553132
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$46897196 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
XM0 2 3 1 4 pfet_03v3 L=2.8e-07 W=2.115e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pmos_1p2$$46898220
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_1p2$$46551084
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sa 1 vss 3 4 qn qp 7 pcb vdd d db se
** N=105 EP=12 IP=47 FDC=27
XM0 1 vss vss vss nfet_03v3 L=2.8e-07 W=1.59e-06 AD=8.866e-13 AS=1.5004e-12 PD=3.93e-06 PS=7.7e-06 NRD=0.0762463 NRS=0.129032 m=1 nf=1 $X=11660 $Y=16585 $D=2
XM1 3 4 1 vss nfet_03v3 L=2.8e-07 W=1.59e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=12780 $Y=16585 $D=2
XM2 4 1 3 vss nfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=1.7732e-12 PD=7.86e-06 PS=7.86e-06 NRD=0.152493 NRS=0.152493 m=1 nf=2 $X=13900 $Y=16585 $D=2
XM3 7 4 vss vss nfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=15170 $Y=8510 $D=2
XM4 1 4 3 vss nfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=1.7732e-12 PD=7.86e-06 PS=7.86e-06 NRD=0.152493 NRS=0.152493 m=1 nf=2 $X=16140 $Y=16585 $D=2
XM5 4 1 3 vss nfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=1.7732e-12 PD=7.86e-06 PS=7.86e-06 NRD=0.152493 NRS=0.152493 m=1 nf=2 $X=18380 $Y=16585 $D=2
XM6 vss 7 qp vss nfet_03v3 L=2.8e-07 W=3.175e-06 AD=1.7706e-12 AS=2.1792e-12 PD=8.37e-06 PS=1.1e-05 NRD=0.343612 NRS=0.422907 m=1 nf=3 $X=17410 $Y=8510 $D=2
XM7 1 4 3 vss nfet_03v3 L=2.8e-07 W=1.59e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=20620 $Y=16585 $D=2
XM8 qn 1 vss vss nfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=20770 $Y=8510 $D=2
XM9 3 se vss vss nfet_03v3 L=2.8e-07 W=1.06e-05 AD=5.9072e-12 AS=6.9296e-12 PD=2.688e-05 PS=3.328e-05 NRD=0.732394 NRS=0.859155 m=1 nf=8 $X=12945 $Y=12550 $D=2
XM10 vss vss 1 vss nfet_03v3 L=2.8e-07 W=1.59e-06 AD=1.5004e-12 AS=8.866e-13 PD=7.7e-06 PS=3.93e-06 NRD=0.129032 NRS=0.0762463 m=1 nf=1 $X=21740 $Y=16585 $D=2
XM11 4 vdd vdd vdd pfet_03v3 L=2.8e-07 W=4.2e-07 AD=2.366e-13 AS=4.004e-13 PD=1.43e-06 PS=2.7e-06 NRD=0.285714 NRS=0.483516 m=1 nf=1 $X=13985 $Y=24010 $D=8
XM12 vdd 1 4 vdd pfet_03v3 L=2.8e-07 W=4.2e-07 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=15105 $Y=24010 $D=8
XM13 d pcb vdd vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=15755 $Y=30660 $D=8
XM14 7 4 vdd vdd pfet_03v3 L=2.8e-07 W=2.115e-06 AD=1.1804e-12 AS=1.589e-12 PD=5.58e-06 PS=8.21e-06 NRD=0.229075 NRS=0.30837 m=1 nf=2 $X=15170 $Y=4385 $D=8
XM15 4 pcb 1 vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=16875 $Y=26330 $D=8
XM16 db pcb d vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=16875 $Y=30660 $D=8
XM17 1 4 vdd vdd pfet_03v3 L=2.8e-07 W=8.45e-07 AD=4.732e-13 AS=4.732e-13 PD=2.86e-06 PS=2.86e-06 NRD=0.571429 NRS=0.571429 m=1 nf=2 $X=16225 $Y=24010 $D=8
XM18 vdd pcb db vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=17995 $Y=30660 $D=8
XM19 4 1 vdd vdd pfet_03v3 L=2.8e-07 W=4.2e-07 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=18465 $Y=24010 $D=8
XM20 qp 7 vdd vdd pfet_03v3 L=2.8e-07 W=2.115e-06 AD=1.1804e-12 AS=1.1804e-12 PD=5.58e-06 PS=5.58e-06 NRD=0.229075 NRS=0.229075 m=1 nf=2 $X=17410 $Y=4385 $D=8
XM21 vdd vdd 4 vdd pfet_03v3 L=2.8e-07 W=4.2e-07 AD=4.004e-13 AS=2.366e-13 PD=2.7e-06 PS=1.43e-06 NRD=0.483516 NRS=0.285714 m=1 nf=1 $X=19585 $Y=24010 $D=8
XM22 qn 1 vdd vdd pfet_03v3 L=2.8e-07 W=2.115e-06 AD=1.1804e-12 AS=1.589e-12 PD=5.58e-06 PS=8.21e-06 NRD=0.229075 NRS=0.30837 m=1 nf=2 $X=19650 $Y=4385 $D=8
X28 db 1 se vdd pmos_1p2$$46897196 $T=12475 26330 0 0 $X=11045 $Y=25620
X29 d 4 se vdd pmos_1p2$$46897196 $T=12475 30660 0 0 $X=11045 $Y=29950
X30 d 4 se vdd pmos_1p2$$46897196 $T=20400 26330 0 0 $X=18970 $Y=25620
X31 db 1 se vdd pmos_1p2$$46897196 $T=20400 30660 0 0 $X=18970 $Y=29950
.ENDS
***************************************
.SUBCKT saout_m2 1 VSS q datain pcb men VDD b[0] bb[0] WEN b[7] bb[7] bb[6] b[6] b[5] bb[5] bb[4] b[4] b[3] bb[3]
+ bb[2] b[2] b[1] bb[1] 54 GWE ypass[7] ypass[6] ypass[5] ypass[4] ypass[3] ypass[2] ypass[1] ypass[0] GWEN 78 79 80 81 82
+ 83 84
** N=135 EP=42 IP=161 FDC=187
*.SEEDPROM
X0 VSS 54 b[0] 74 bb[0] 77 pcb VDD ypass[0] 78 bb[7] b[7] 79 bb[6] b[6] 80 bb[5] b[5] 81 bb[4]
+ b[4] 82 bb[3] b[3] 83 bb[2] b[2] 84 bb[1] b[1] ypass[7] ypass[6] ypass[5] ypass[4] ypass[3] ypass[2] ypass[1]
+ mux821 $T=2765 83345 0 0 $X=-1345 $Y=83340
X1 VSS 1 86 89 90 87 92 96 91 97 93 94 95 men VDD WEN GWEN 85 88 wen_wm1 $T=1610 -16845 0 0 $X=100 $Y=-17385
X2 VSS 98 pcb 72 103 104 105 106 108 111 112 100 99 101 75 102 73 107 109 110
+ 76 VDD men
+ sacntl_2 $T=3160 150 0 0 $X=425 $Y=30
X3 q VSS 113 115 116 118 117 114 120 VDD GWE 76 134 135 119 outbuf_oe $T=3160 27580 0 0 $X=500 $Y=25785
X4 VSS 121 124 129 74 77 126 122 125 127 128 123 VDD datain men 1 din $T=1615 39060 0 0 $X=500 $Y=38775
X5 130 VSS 132 131 135 134 133 pcb VDD 74 77 76 sa $T=3160 43075 0 0 $X=1375 $Y=42095
.ENDS
***************************************
.SUBCKT 018SRAM_cell1_dummy 1 2 3 4 5 7
** N=9 EP=6 IP=0 FDC=4
*.SEEDPROM
XM0 1 7 2 3 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=180 $Y=260 $D=2
XM1 3 5 1 3 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=1710 $D=2
XM2 5 1 3 3 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=1710 $D=2
XM3 5 7 4 3 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=2220 $Y=260 $D=2
.ENDS
***************************************
.SUBCKT ICV_7 1 3 4 5 6 7 8 9 10 11
** N=15 EP=10 IP=18 FDC=8
*.SEEDPROM
X0 5 4 1 6 7 3 018SRAM_cell1_dummy $T=-3000 0 0 0 $X=-3340 $Y=-340
X1 9 8 1 10 11 3 018SRAM_cell1_dummy $T=0 0 0 0 $X=-340 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_8 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19
** N=27 EP=18 IP=30 FDC=16
*.SEEDPROM
X0 1 3 4 5 6 7 8 9 10 11 ICV_7 $T=-6000 0 0 0 $X=-9340 $Y=-340
X1 1 3 12 13 14 15 16 17 18 19 ICV_7 $T=0 0 0 0 $X=-3340 $Y=-340
.ENDS
***************************************
.SUBCKT 018SRAM_strap1
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
** N=30 EP=18 IP=33 FDC=16
*.SEEDPROM
X0 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 ICV_8 $T=-3000 0 0 0 $X=-12340 $Y=-340
.ENDS
***************************************
.SUBCKT 018SRAM_cell1
** N=8 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT 018SRAM_cell1_2x 1 2 3 5 6 7 8 9 10
** N=12 EP=9 IP=16 FDC=8
*.SEEDPROM
XM0 1 5 7 3 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=180 $Y=3470 $D=2
XM1 9 6 1 3 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=180 $Y=4760 $D=2
XM2 3 8 7 3 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=1840 $D=2
XM3 3 10 9 3 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=6210 $D=2
XM4 8 7 3 3 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=1840 $D=2
XM5 10 9 3 3 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=6210 $D=2
XM6 2 5 8 3 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=2220 $Y=3470 $D=2
XM7 10 6 2 3 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=2220 $Y=4760 $D=2
.ENDS
***************************************
.SUBCKT ICV_11 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
** N=16 EP=15 IP=24 FDC=16
*.SEEDPROM
X0 5 6 2 3 4 9 11 10 12 018SRAM_cell1_2x $T=0 0 0 0 $X=-340 $Y=-340
X1 7 8 2 3 4 13 15 14 16 018SRAM_cell1_2x $T=3000 0 0 0 $X=2660 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_12 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=26 EP=18 IP=32 FDC=40
*.SEEDPROM
XM0 1 20 19 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=8060 $D=8
XM1 1 24 23 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=9340 $D=8
XM2 20 19 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=8060 $D=8
XM3 24 23 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=9340 $D=8
XM4 1 22 21 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=8060 $D=8
XM5 1 26 25 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=9340 $D=8
XM6 22 21 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=8060 $D=8
XM7 26 25 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=9340 $D=8
X8 2 3 4 7 8 9 10 11 19 12 20 13 21 14 22 ICV_11 $T=0 0 0 0 $X=-340 $Y=-340
X9 2 5 6 7 8 9 10 23 15 24 16 25 17 26 18 ICV_11 $T=0 9000 0 0 $X=-340 $Y=8660
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
** N=30 EP=30 IP=36 FDC=80
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 15 16 17 18 19 20 21 22 ICV_12 $T=0 0 0 0 $X=-340 $Y=-340
X1 1 2 3 4 5 6 11 12 13 14 23 24 25 26 27 28 29 30 ICV_12 $T=6000 0 0 0 $X=5660 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_14 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34
** N=50 EP=34 IP=60 FDC=176
*.SEEDPROM
XM0 1 36 35 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=17060 $D=8
XM1 1 44 43 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=18340 $D=8
XM2 36 35 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=17060 $D=8
XM3 44 43 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=18340 $D=8
XM4 1 38 37 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=17060 $D=8
XM5 1 46 45 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=18340 $D=8
XM6 38 37 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=17060 $D=8
XM7 46 45 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=18340 $D=8
XM8 1 40 39 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=6630 $Y=17060 $D=8
XM9 1 48 47 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=6630 $Y=18340 $D=8
XM10 40 39 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=7770 $Y=17060 $D=8
XM11 48 47 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=7770 $Y=18340 $D=8
XM12 1 42 41 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=9630 $Y=17060 $D=8
XM13 1 50 49 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=9630 $Y=18340 $D=8
XM14 42 41 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=10770 $Y=17060 $D=8
XM15 50 49 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=10770 $Y=18340 $D=8
X16 1 2 3 4 5 6 11 12 13 14 15 16 17 18 19 20 21 22 35 36
+ 37 38 23 24 25 26 39 40 41 42
+ ICV_13 $T=0 0 0 0 $X=-340 $Y=-340
X17 1 2 7 8 9 10 11 12 13 14 15 16 17 18 43 44 45 46 27 28
+ 29 30 47 48 49 50 31 32 33 34
+ ICV_13 $T=0 18000 0 0 $X=-340 $Y=17660
.ENDS
***************************************
.SUBCKT 018SRAM_strap1_2x
** N=10 EP=0 IP=12 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=15 EP=0 IP=20 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16
** N=19 EP=0 IP=24 FDC=0
.ENDS
***************************************
.SUBCKT ICV_25 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 27 28 29 30 31 32 33 34 35 36 37 38 39 40
** N=40 EP=34 IP=50 FDC=176
*.SEEDPROM
X0 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ ICV_14 $T=0 -4500 1 180 $X=-12340 $Y=-4840
.ENDS
***************************************
.SUBCKT ICV_26 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 27 28 29 30 31 32 36 37 38 39 40 41 42 43 44 45 46 47 48 49
+ 50 51
** N=67 EP=42 IP=80 FDC=368
*.SEEDPROM
XM0 7 58 59 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-11370 $Y=30560 $D=8
XM1 7 66 67 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-11370 $Y=31840 $D=8
XM2 58 59 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-10230 $Y=30560 $D=8
XM3 66 67 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-10230 $Y=31840 $D=8
XM4 7 56 57 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-8370 $Y=30560 $D=8
XM5 7 64 65 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-8370 $Y=31840 $D=8
XM6 56 57 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-7230 $Y=30560 $D=8
XM7 64 65 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-7230 $Y=31840 $D=8
XM8 7 54 55 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-5370 $Y=30560 $D=8
XM9 7 62 63 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-5370 $Y=31840 $D=8
XM10 54 55 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-4230 $Y=30560 $D=8
XM11 62 63 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-4230 $Y=31840 $D=8
XM12 7 52 53 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=30560 $D=8
XM13 7 60 61 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=31840 $D=8
XM14 52 53 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=30560 $D=8
XM15 60 61 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=31840 $D=8
X16 7 8 9 10 11 12 13 14 15 16 32 31 30 29 28 27 26 25 36 37
+ 38 39 40 41 42 43 52 53 54 55 56 57 58 59
+ ICV_25 $T=0 0 0 0 $X=-12340 $Y=-4840
X17 7 8 17 18 19 20 21 22 23 24 32 31 30 29 28 27 26 25 60 61
+ 62 63 64 65 66 67 44 45 46 47 48 49 50 51
+ ICV_25 $T=0 36000 0 0 $X=-12340 $Y=31160
.ENDS
***************************************
.SUBCKT ICV_27 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46
+ 47 48 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67
** N=83 EP=58 IP=96 FDC=752
*.SEEDPROM
XM0 7 74 75 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-11370 $Y=66560 $D=8
XM1 7 82 83 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-11370 $Y=67840 $D=8
XM2 74 75 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-10230 $Y=66560 $D=8
XM3 82 83 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-10230 $Y=67840 $D=8
XM4 7 72 73 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-8370 $Y=66560 $D=8
XM5 7 80 81 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-8370 $Y=67840 $D=8
XM6 72 73 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-7230 $Y=66560 $D=8
XM7 80 81 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-7230 $Y=67840 $D=8
XM8 7 70 71 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-5370 $Y=66560 $D=8
XM9 7 78 79 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-5370 $Y=67840 $D=8
XM10 70 71 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-4230 $Y=66560 $D=8
XM11 78 79 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-4230 $Y=67840 $D=8
XM12 7 68 69 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=66560 $D=8
XM13 7 76 77 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=67840 $D=8
XM14 68 69 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=66560 $D=8
XM15 76 77 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=67840 $D=8
X16 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 41 42
+ 43 44 45 46 47 48 52 53 54 55 56 57 58 59 68 69 70 71 72 73
+ 74 75
+ ICV_26 $T=0 0 0 0 $X=-12340 $Y=-4840
X17 7 8 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 76 77 78 79 80 81 82 83 60 61 62 63 64 65
+ 66 67
+ ICV_26 $T=0 72000 0 0 $X=-12340 $Y=67160
.ENDS
***************************************
.SUBCKT ICV_10 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35 36 37 38
** N=54 EP=34 IP=57 FDC=32
*.SEEDPROM
X0 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 ICV_8 $T=-15000 0 0 0 $X=-24340 $Y=-340
X1 4 6 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 ICV_9 $T=0 0 0 0 $X=-12340 $Y=-340
.ENDS
***************************************
.SUBCKT dcap_103_novia
** N=2 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_5
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_6
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_17 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 27 28 29 30 31 32 33 34 35 36 37 38 39 40
** N=40 EP=34 IP=50 FDC=176
*.SEEDPROM
X0 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ ICV_14 $T=0 0 0 0 $X=-340 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_18 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
** N=16 EP=15 IP=24 FDC=16
*.SEEDPROM
X0 5 6 2 3 4 9 11 10 12 018SRAM_cell1_2x $T=-3000 0 0 0 $X=-3340 $Y=-340
X1 7 8 2 3 4 13 15 14 16 018SRAM_cell1_2x $T=0 0 0 0 $X=-340 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_19 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=26 EP=18 IP=32 FDC=40
*.SEEDPROM
XM0 1 20 19 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=8060 $D=8
XM1 1 24 23 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=9340 $D=8
XM2 20 19 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=8060 $D=8
XM3 24 23 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=9340 $D=8
XM4 1 22 21 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=8060 $D=8
XM5 1 26 25 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=9340 $D=8
XM6 22 21 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=8060 $D=8
XM7 26 25 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=9340 $D=8
X8 2 3 4 7 8 9 10 11 19 12 20 13 21 14 22 ICV_18 $T=0 0 0 0 $X=-3340 $Y=-340
X9 2 5 6 7 8 9 10 23 15 24 16 25 17 26 18 ICV_18 $T=0 9000 0 0 $X=-3340 $Y=8660
.ENDS
***************************************
.SUBCKT ICV_20 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
** N=30 EP=30 IP=36 FDC=80
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 15 16 17 18 19 20 21 22 ICV_19 $T=-6000 0 0 0 $X=-9340 $Y=-340
X1 1 2 3 4 5 6 11 12 13 14 23 24 25 26 27 28 29 30 ICV_19 $T=0 0 0 0 $X=-3340 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_21 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34
** N=50 EP=34 IP=60 FDC=176
*.SEEDPROM
XM0 1 36 35 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-8370 $Y=17060 $D=8
XM1 1 44 43 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-8370 $Y=18340 $D=8
XM2 36 35 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-7230 $Y=17060 $D=8
XM3 44 43 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-7230 $Y=18340 $D=8
XM4 1 38 37 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-5370 $Y=17060 $D=8
XM5 1 46 45 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-5370 $Y=18340 $D=8
XM6 38 37 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-4230 $Y=17060 $D=8
XM7 46 45 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-4230 $Y=18340 $D=8
XM8 1 40 39 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=17060 $D=8
XM9 1 48 47 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=18340 $D=8
XM10 40 39 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=17060 $D=8
XM11 48 47 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=18340 $D=8
XM12 1 42 41 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=17060 $D=8
XM13 1 50 49 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=18340 $D=8
XM14 42 41 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=17060 $D=8
XM15 50 49 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=18340 $D=8
X16 1 2 3 4 5 6 11 12 13 14 15 16 17 18 19 20 21 22 35 36
+ 37 38 23 24 25 26 39 40 41 42
+ ICV_20 $T=0 0 0 0 $X=-9340 $Y=-340
X17 1 2 7 8 9 10 11 12 13 14 15 16 17 18 43 44 45 46 27 28
+ 29 30 47 48 49 50 31 32 33 34
+ ICV_20 $T=0 18000 0 0 $X=-9340 $Y=17660
.ENDS
***************************************
.SUBCKT ICV_22 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58
** N=58 EP=58 IP=68 FDC=352
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 27 28
+ 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ ICV_21 $T=-12000 0 0 0 $X=-21340 $Y=-340
X1 1 2 3 4 5 6 7 8 9 10 19 20 21 22 23 24 25 26 43 44
+ 45 46 47 48 49 50 51 52 53 54 55 56 57 58
+ ICV_21 $T=0 0 0 0 $X=-9340 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_23 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46
+ 47 48 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69
+ 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89
+ 90 91 92 93 94 95 96 97 98 99
** N=147 EP=90 IP=196 FDC=1104
*.SEEDPROM
XM0 7 101 100 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=35060 $D=8
XM1 7 109 108 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=36340 $D=8
XM2 101 100 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=35060 $D=8
XM3 109 108 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=36340 $D=8
XM4 7 103 102 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=35060 $D=8
XM5 7 111 110 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=36340 $D=8
XM6 103 102 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=35060 $D=8
XM7 111 110 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=36340 $D=8
XM8 7 105 104 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=6630 $Y=35060 $D=8
XM9 7 113 112 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=6630 $Y=36340 $D=8
XM10 105 104 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=7770 $Y=35060 $D=8
XM11 113 112 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=7770 $Y=36340 $D=8
XM12 7 107 106 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=9630 $Y=35060 $D=8
XM13 7 115 114 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=9630 $Y=36340 $D=8
XM14 107 106 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=10770 $Y=35060 $D=8
XM15 115 114 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=10770 $Y=36340 $D=8
XM16 7 130 131 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15630 $Y=35060 $D=8
XM17 7 146 147 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15630 $Y=36340 $D=8
XM18 130 131 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16770 $Y=35060 $D=8
XM19 146 147 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16770 $Y=36340 $D=8
XM20 7 128 129 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18630 $Y=35060 $D=8
XM21 7 144 145 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18630 $Y=36340 $D=8
XM22 128 129 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19770 $Y=35060 $D=8
XM23 144 145 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19770 $Y=36340 $D=8
XM24 7 126 127 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21630 $Y=35060 $D=8
XM25 7 142 143 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21630 $Y=36340 $D=8
XM26 126 127 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22770 $Y=35060 $D=8
XM27 142 143 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22770 $Y=36340 $D=8
XM28 7 124 125 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24630 $Y=35060 $D=8
XM29 7 140 141 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24630 $Y=36340 $D=8
XM30 124 125 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25770 $Y=35060 $D=8
XM31 140 141 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25770 $Y=36340 $D=8
XM32 7 122 123 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27630 $Y=35060 $D=8
XM33 7 138 139 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27630 $Y=36340 $D=8
XM34 122 123 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28770 $Y=35060 $D=8
XM35 138 139 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28770 $Y=36340 $D=8
XM36 7 120 121 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30630 $Y=35060 $D=8
XM37 7 136 137 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30630 $Y=36340 $D=8
XM38 120 121 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31770 $Y=35060 $D=8
XM39 136 137 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31770 $Y=36340 $D=8
XM40 7 118 119 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33630 $Y=35060 $D=8
XM41 7 134 135 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33630 $Y=36340 $D=8
XM42 118 119 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34770 $Y=35060 $D=8
XM43 134 135 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34770 $Y=36340 $D=8
XM44 7 116 117 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=36630 $Y=35060 $D=8
XM45 7 132 133 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=36630 $Y=36340 $D=8
XM46 116 117 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=37770 $Y=35060 $D=8
XM47 132 133 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=37770 $Y=36340 $D=8
X48 7 8 9 10 11 12 13 14 15 16 25 26 27 28 29 30 31 32 52 53
+ 54 55 56 57 58 59 100 101 102 103 104 105 106 107
+ ICV_17 $T=0 0 0 0 $X=-340 $Y=-340
X49 7 8 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 108 109
+ 110 111 112 113 114 115 60 61 62 63 64 65 66 67
+ ICV_17 $T=0 36000 0 0 $X=-340 $Y=35660
X50 7 8 9 10 11 12 13 14 15 16 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 68 69 70 71 72 73 74 75 116 117 118 119 120 121
+ 122 123 76 77 78 79 80 81 82 83 124 125 126 127 128 129 130 131
+ ICV_22 $T=18000 0 1 180 $X=14660 $Y=-340
X51 7 8 17 18 19 20 21 22 23 24 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 132 133 134 135 136 137 138 139 84 85 86 87 88 89
+ 90 91 140 141 142 143 144 145 146 147 92 93 94 95 96 97 98 99
+ ICV_22 $T=18000 36000 1 180 $X=14660 $Y=35660
.ENDS
***************************************
.SUBCKT ICV_24 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46
+ 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 68 69
+ 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89
+ 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109
+ 110 111 112 113 114 115
** N=163 EP=106 IP=192 FDC=2256
*.SEEDPROM
XM0 7 117 116 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=71060 $D=8
XM1 7 141 140 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=72340 $D=8
XM2 117 116 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=71060 $D=8
XM3 141 140 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=72340 $D=8
XM4 7 119 118 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=71060 $D=8
XM5 7 143 142 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=72340 $D=8
XM6 119 118 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=71060 $D=8
XM7 143 142 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=72340 $D=8
XM8 7 121 120 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=6630 $Y=71060 $D=8
XM9 7 145 144 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=6630 $Y=72340 $D=8
XM10 121 120 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=7770 $Y=71060 $D=8
XM11 145 144 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=7770 $Y=72340 $D=8
XM12 7 123 122 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=9630 $Y=71060 $D=8
XM13 7 147 146 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=9630 $Y=72340 $D=8
XM14 123 122 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=10770 $Y=71060 $D=8
XM15 147 146 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=10770 $Y=72340 $D=8
XM16 7 138 139 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15630 $Y=71060 $D=8
XM17 7 162 163 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15630 $Y=72340 $D=8
XM18 138 139 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16770 $Y=71060 $D=8
XM19 162 163 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16770 $Y=72340 $D=8
XM20 7 136 137 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18630 $Y=71060 $D=8
XM21 7 160 161 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18630 $Y=72340 $D=8
XM22 136 137 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19770 $Y=71060 $D=8
XM23 160 161 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19770 $Y=72340 $D=8
XM24 7 134 135 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21630 $Y=71060 $D=8
XM25 7 158 159 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21630 $Y=72340 $D=8
XM26 134 135 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22770 $Y=71060 $D=8
XM27 158 159 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22770 $Y=72340 $D=8
XM28 7 132 133 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24630 $Y=71060 $D=8
XM29 7 156 157 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24630 $Y=72340 $D=8
XM30 132 133 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25770 $Y=71060 $D=8
XM31 156 157 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25770 $Y=72340 $D=8
XM32 7 130 131 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27630 $Y=71060 $D=8
XM33 7 154 155 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27630 $Y=72340 $D=8
XM34 130 131 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28770 $Y=71060 $D=8
XM35 154 155 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28770 $Y=72340 $D=8
XM36 7 128 129 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30630 $Y=71060 $D=8
XM37 7 152 153 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30630 $Y=72340 $D=8
XM38 128 129 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31770 $Y=71060 $D=8
XM39 152 153 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31770 $Y=72340 $D=8
XM40 7 126 127 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33630 $Y=71060 $D=8
XM41 7 150 151 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33630 $Y=72340 $D=8
XM42 126 127 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34770 $Y=71060 $D=8
XM43 150 151 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34770 $Y=72340 $D=8
XM44 7 124 125 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=36630 $Y=71060 $D=8
XM45 7 148 149 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=36630 $Y=72340 $D=8
XM46 124 125 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=37770 $Y=71060 $D=8
XM47 148 149 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=37770 $Y=72340 $D=8
X48 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 41 42
+ 43 44 45 46 47 48 64 63 62 61 60 59 58 57 56 55 54 53 52 51
+ 50 49 68 69 70 71 72 73 74 75 116 117 118 119 120 121 122 123 76 77
+ 78 79 80 81 82 83 84 85 86 87 88 89 90 91 124 125 126 127 128 129
+ 130 131 132 133 134 135 136 137 138 139
+ ICV_23 $T=0 0 0 0 $X=-340 $Y=-340
X49 7 8 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 64 63 62 61 60 59 58 57 56 55 54 53 52 51
+ 50 49 140 141 142 143 144 145 146 147 92 93 94 95 96 97 98 99 148 149
+ 150 151 152 153 154 155 156 157 158 159 160 161 162 163 100 101 102 103 104 105
+ 106 107 108 109 110 111 112 113 114 115
+ ICV_23 $T=0 72000 0 0 $X=-340 $Y=71660
.ENDS
***************************************
.SUBCKT saout_R_m2 1 vss q pcb datain men vdd b[7] bb[7] WEN b[0] bb[0] bb[1] b[1] b[2] bb[2] bb[3] b[3] b[4] bb[4]
+ bb[5] b[5] b[6] bb[6] 54 GWE ypass[0] ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] GWEN 74 75 76 77 78
+ 79 80
** N=131 EP=42 IP=161 FDC=187
*.SEEDPROM
X0 vss 54 b[7] 70 bb[7] 73 pcb vdd ypass[7] 74 bb[0] b[0] 75 bb[1] b[1] 76 bb[2] b[2] 77 bb[3]
+ b[3] 78 bb[4] b[4] 79 bb[5] b[5] 80 bb[6] b[6] ypass[0] ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6]
+ mux821 $T=2765 83310 0 0 $X=-1345 $Y=83305
X1 vss 1 82 85 86 83 88 92 87 93 89 90 91 men vdd WEN GWEN 81 84 wen_wm1 $T=1610 -16880 0 0 $X=100 $Y=-17420
X2 vss 94 pcb 68 99 100 101 102 104 107 108 96 95 97 71 98 69 103 105 106
+ 72 vdd men
+ sacntl_2 $T=3160 115 0 0 $X=425 $Y=-5
X3 q vss 109 111 112 114 113 110 116 vdd GWE 72 130 131 115 outbuf_oe $T=3160 27545 0 0 $X=500 $Y=25750
X4 vss 117 120 125 70 73 122 118 121 123 124 119 vdd datain men 1 din $T=1615 39025 0 0 $X=500 $Y=38740
X5 126 vss 128 127 131 130 129 pcb vdd 70 73 72 sa $T=3160 43040 0 0 $X=1375 $Y=42060
.ENDS
***************************************
.SUBCKT 018SRAM_strap1_bndry
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT 018SRAM_strap1_2x_bndry
** N=10 EP=0 IP=12 FDC=0
.ENDS
***************************************
.SUBCKT ICV_38
** N=15 EP=0 IP=20 FDC=0
.ENDS
***************************************
.SUBCKT 018SRAM_cell1_cutPC
** N=7 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_39 1 2 4 7 8 9 10
** N=10 EP=7 IP=14 FDC=8
*.SEEDPROM
XM0 1 4 7 4 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=180 $Y=-1030 $D=2
XM1 9 4 1 4 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=180 $Y=260 $D=2
XM2 4 8 7 4 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=-2660 $D=2
XM3 4 10 9 4 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=1710 $D=2
XM4 8 7 4 4 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=-2660 $D=2
XM5 10 9 4 4 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=1710 $D=2
XM6 2 4 8 4 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=2220 $Y=-1030 $D=2
XM7 10 4 2 4 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=2220 $Y=260 $D=2
.ENDS
***************************************
.SUBCKT ICV_40 1 2 7 8 9 10 11 12
** N=16 EP=8 IP=20 FDC=20
*.SEEDPROM
XM0 1 14 13 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=-5440 $D=8
XM1 1 16 15 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=-4160 $D=8
XM2 14 13 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=-5440 $D=8
XM3 16 15 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=-4160 $D=8
X4 7 8 2 9 10 13 14 ICV_39 $T=0 -9000 0 0 $X=-340 $Y=-13840
X5 7 8 2 15 16 11 12 ICV_39 $T=0 0 0 0 $X=-340 $Y=-4840
.ENDS
***************************************
.SUBCKT ICV_41 7 8 17 18 22 23 24 25
** N=29 EP=8 IP=48 FDC=44
*.SEEDPROM
XM0 7 26 27 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=12560 $D=8
XM1 7 28 29 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=13840 $D=8
XM2 26 27 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=12560 $D=8
XM3 28 29 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=13840 $D=8
X6 7 8 17 18 26 27 22 23 ICV_40 $T=6000 0 0 180 $X=2660 $Y=-4840
X7 7 8 17 18 24 25 28 29 ICV_40 $T=6000 18000 0 180 $X=2660 $Y=13160
.ENDS
***************************************
.SUBCKT pfet_03v3_I07
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT M1_POLY2_I01
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nfet_03v3_I03
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2_01_R270 1 2 3
** N=3 EP=3 IP=0 FDC=1
XM0 2 3 1 1 pfet_03v3 L=2.8e-07 W=5.13e-06 AD=2.86e-12 AS=4.84e-12 PD=1.204e-05 PS=2.376e-05 NRD=0.0945455 NRS=0.16 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pfet_03v3_I05
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT xdec 1 2 men 6 vss 8 28 vdd
** N=104 EP=8 IP=41 FDC=6
*.SEEDPROM
XM0 2 6 men vss nfet_03v3 L=2.8e-07 W=3.08e-06 AD=2.904e-12 AS=1.716e-12 PD=1.496e-05 PS=7.64e-06 NRD=0.266667 NRS=0.157576 m=1 nf=2 $X=37460 $Y=965 $D=2
XM1 vss 8 6 vss nfet_03v3 L=2.8e-07 W=3.05e-07 AD=2.904e-13 AS=2.904e-13 PD=2.2e-06 PS=2.2e-06 NRD=0.666667 NRS=0.666667 m=1 nf=1 $X=45970 $Y=965 $D=2
XM2 2 8 men vdd pfet_03v3 L=2.8e-07 W=3.08e-06 AD=2.904e-12 AS=1.716e-12 PD=1.496e-05 PS=7.64e-06 NRD=0.266667 NRS=0.157576 m=1 nf=2 $X=32185 $Y=965 $D=8
XM3 vdd 8 6 vdd pfet_03v3 L=2.8e-07 W=7.4e-07 AD=6.996e-13 AS=6.996e-13 PD=4.06e-06 PS=4.06e-06 NRD=0.27673 NRS=0.27673 m=1 nf=1 $X=43020 $Y=965 $D=8
X12 vdd 1 2 pmos_1p2_01_R270 $T=29780 1120 0 90 $X=23605 $Y=-360
X13 vdd 28 2 pmos_1p2_01_R270 $T=91805 1120 1 90 $X=91120 $Y=-360
.ENDS
***************************************
.SUBCKT xdec8 vss xc xb xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] vdd 102 men 104 LWL[1] RWL[1] LWL[2] RWL[2] LWL[3] RWL[3] LWL[4]
+ RWL[4] LWL[5] RWL[5] LWL[6] RWL[6] 120 121 270 273 316 319
** N=335 EP=31 IP=616 FDC=126
*.SEEDPROM
XM0 vss 275 274 vss nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=16340 $Y=5740 $D=2
XM1 vss 274 LWL[1] vss nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=7020 $D=2
XM2 vss 281 LWL[2] vss nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=9260 $D=2
XM3 281 282 vss vss nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=16340 $Y=11660 $D=2
XM4 vss 289 288 vss nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=16340 $Y=14740 $D=2
XM5 vss 288 LWL[3] vss nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=16020 $D=2
XM6 vss 295 LWL[4] vss nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=18260 $D=2
XM7 295 296 vss vss nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=16340 $Y=20660 $D=2
XM8 vss 303 302 vss nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=16340 $Y=23740 $D=2
XM9 vss 302 LWL[5] vss nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=25020 $D=2
XM10 vss 309 LWL[6] vss nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=27260 $D=2
XM11 309 310 vss vss nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=16340 $Y=29660 $D=2
XM12 vss 277 275 vss nfet_03v3 L=2.8e-07 W=1.025e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=46620 $Y=8140 $D=2
XM13 282 284 vss vss nfet_03v3 L=2.8e-07 W=1.025e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=46620 $Y=9260 $D=2
XM14 vss 291 289 vss nfet_03v3 L=2.8e-07 W=1.025e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=46620 $Y=17140 $D=2
XM15 296 298 vss vss nfet_03v3 L=2.8e-07 W=1.025e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=46620 $Y=18260 $D=2
XM16 vss 305 303 vss nfet_03v3 L=2.8e-07 W=1.025e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=46620 $Y=26140 $D=2
XM17 310 312 vss vss nfet_03v3 L=2.8e-07 W=1.025e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=46620 $Y=27260 $D=2
XM18 324 xa[1] 277 vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=66460 $Y=5900 $D=2
XM19 325 xb 324 vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=66460 $Y=7020 $D=2
XM20 vss xc 325 vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=66460 $Y=8085 $D=2
XM21 327 xc vss vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=66460 $Y=9315 $D=2
XM22 326 xb 327 vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=66460 $Y=10380 $D=2
XM23 284 xa[2] 326 vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=66460 $Y=11500 $D=2
XM24 328 xa[3] 291 vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=66460 $Y=14900 $D=2
XM25 329 xb 328 vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=66460 $Y=16020 $D=2
XM26 vss xc 329 vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=66460 $Y=17085 $D=2
XM27 331 xc vss vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=66460 $Y=18315 $D=2
XM28 330 xb 331 vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=66460 $Y=19380 $D=2
XM29 298 xa[4] 330 vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=66460 $Y=20500 $D=2
XM30 332 xa[5] 305 vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=66460 $Y=23900 $D=2
XM31 333 xb 332 vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=66460 $Y=25020 $D=2
XM32 vss xc 333 vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=66460 $Y=26085 $D=2
XM33 335 xc vss vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=66460 $Y=27315 $D=2
XM34 334 xb 335 vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=66460 $Y=28380 $D=2
XM35 312 xa[6] 334 vss nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=66460 $Y=29500 $D=2
XM36 vss 275 280 vss nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=100255 $Y=5740 $D=2
XM37 vss 280 RWL[1] vss nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=7020 $D=2
XM38 vss 287 RWL[2] vss nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=9260 $D=2
XM39 287 282 vss vss nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=100255 $Y=11660 $D=2
XM40 vss 289 294 vss nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=100255 $Y=14740 $D=2
XM41 vss 294 RWL[3] vss nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=16020 $D=2
XM42 vss 301 RWL[4] vss nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=18260 $D=2
XM43 301 296 vss vss nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=100255 $Y=20660 $D=2
XM44 vss 303 308 vss nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=100255 $Y=23740 $D=2
XM45 vss 308 RWL[5] vss nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=25020 $D=2
XM46 vss 315 RWL[6] vss nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=27260 $D=2
XM47 315 310 vss vss nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=100255 $Y=29660 $D=2
XM48 LWL[1] 274 vdd vdd pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=4665 $Y=5900 $D=8
XM49 vdd 281 LWL[2] vdd pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=4665 $Y=9260 $D=8
XM50 LWL[3] 288 vdd vdd pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=4665 $Y=14900 $D=8
XM51 vdd 295 LWL[4] vdd pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=4665 $Y=18260 $D=8
XM52 LWL[5] 302 vdd vdd pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=4665 $Y=23900 $D=8
XM53 vdd 309 LWL[6] vdd pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=4665 $Y=27260 $D=8
XM54 vdd xa[1] 277 vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=71980 $Y=5900 $D=8
XM55 277 xb vdd vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=7020 $D=8
XM56 vdd xc 277 vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=8140 $D=8
XM57 284 xc vdd vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=9260 $D=8
XM58 vdd xb 284 vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=10380 $D=8
XM59 284 xa[2] vdd vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=71980 $Y=11500 $D=8
XM60 vdd xa[3] 291 vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=71980 $Y=14900 $D=8
XM61 291 xb vdd vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=16020 $D=8
XM62 vdd xc 291 vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=17140 $D=8
XM63 298 xc vdd vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=18260 $D=8
XM64 vdd xb 298 vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=19380 $D=8
XM65 298 xa[4] vdd vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=71980 $Y=20500 $D=8
XM66 vdd xa[5] 305 vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=71980 $Y=23900 $D=8
XM67 305 xb vdd vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=25020 $D=8
XM68 vdd xc 305 vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=26140 $D=8
XM69 312 xc vdd vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=27260 $D=8
XM70 vdd xb 312 vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=28380 $D=8
XM71 312 xa[6] vdd vdd pfet_03v3 L=2.8e-07 W=1.22e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=71980 $Y=29500 $D=8
XM72 RWL[1] 280 vdd vdd pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=106930 $Y=5900 $D=8
XM73 vdd 287 RWL[2] vdd pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=106930 $Y=9260 $D=8
XM74 RWL[3] 294 vdd vdd pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=106930 $Y=14900 $D=8
XM75 vdd 301 RWL[4] vdd pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=106930 $Y=18260 $D=8
XM76 RWL[5] 308 vdd vdd pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=106930 $Y=23900 $D=8
XM77 vdd 315 RWL[6] vdd pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=106930 $Y=27260 $D=8
X78 270 102 men 271 vss 104 273 vdd xdec $T=5 4500 1 0 $X=0 $Y=-1140
X79 274 275 men 276 vss 277 280 vdd xdec $T=5 4500 0 0 $X=0 $Y=3385
X80 281 282 men 283 vss 284 287 vdd xdec $T=5 13500 1 0 $X=0 $Y=7860
X81 288 289 men 290 vss 291 294 vdd xdec $T=5 13500 0 0 $X=0 $Y=12385
X82 295 296 men 297 vss 298 301 vdd xdec $T=5 22500 1 0 $X=0 $Y=16860
X83 302 303 men 304 vss 305 308 vdd xdec $T=5 22500 0 0 $X=0 $Y=21385
X84 309 310 men 311 vss 312 315 vdd xdec $T=5 31500 1 0 $X=0 $Y=25860
X85 316 120 men 317 vss 121 319 vdd xdec $T=5 31500 0 0 $X=0 $Y=30385
.ENDS
***************************************
.SUBCKT pmoscap_R270
** N=26 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_35
** N=6 EP=0 IP=8 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_36
** N=10 EP=0 IP=12 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_37 1 50 51 52 54 55 56 57 58 59 104 105 106 107 108 109 112 113 114 115
+ 116 117 119 126 127 128 129 130 131 132 133
** N=137 EP=31 IP=157 FDC=126
*.SEEDPROM
X0 1 51 52 59 58 57 56 55 54 50 126 119 127 104 112 105 113 106 114 107
+ 115 108 116 109 117 128 129 130 131 132 133
+ xdec8 $T=9750 2385 1 270 $X=-27390 $Y=-118710
.ENDS
***************************************
.SUBCKT pmoscap_L1_W2_R270
** N=13 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT M1_PSUB_I03
** N=2001 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pmos_1p2$$47513644
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_03v3_I21
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_1p2$$47641644
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pfet_03v3_I12
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT xpredec0_xa 2 3 13 29 30
** N=40 EP=5 IP=40 FDC=4
*.SEEDPROM
XM0 40 29 2 3 nfet_03v3 L=2.8e-07 W=5.715e-06 AD=3.185e-12 AS=7.2275e-12 PD=1.277e-05 PS=2.568e-05 NRD=0.0212245 NRS=0.0481633 m=1 nf=1 $X=3255 $Y=2430 $D=2
XM1 3 30 40 3 nfet_03v3 L=2.8e-07 W=5.715e-06 AD=7.28875e-12 AS=3.185e-12 PD=2.569e-05 PS=1.277e-05 NRD=0.0485714 NRS=0.0212245 m=1 nf=1 $X=4375 $Y=2430 $D=2
XM2 2 29 13 13 pfet_03v3 L=2.8e-07 W=7.09e-06 AD=3.952e-12 AS=6.688e-12 PD=1.572e-05 PS=3.128e-05 NRD=0.0171053 NRS=0.0289474 m=1 nf=1 $X=3255 $Y=19540 $D=8
XM3 13 30 2 13 pfet_03v3 L=2.8e-07 W=7.09e-06 AD=6.688e-12 AS=3.952e-12 PD=3.128e-05 PS=1.572e-05 NRD=0.0289474 NRS=0.0171053 m=1 nf=1 $X=4375 $Y=19540 $D=8
.ENDS
***************************************
.SUBCKT pmos_1p2_161 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
XM0 2 3 1 4 pfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT alatch vss ab a vdd enb en
** N=16 EP=6 IP=24 FDC=8
XM0 ab 12 vss vss nfet_03v3 L=2.8e-07 W=1.695e-06 AD=9.464e-13 AS=1.6016e-12 PD=4.68e-06 PS=9.04e-06 NRD=0.285714 NRS=0.483516 m=1 nf=2 $X=2590 $Y=1475 $D=2
XM1 vss ab 11 vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=3710 $Y=12935 $D=2
XM2 a en 12 vss nfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=6280 $Y=1020 $D=2
XM3 11 enb 12 vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=6280 $Y=12935 $D=2
XM4 ab 12 vdd vdd pfet_03v3 L=2.8e-07 W=4.235e-06 AD=2.3608e-12 AS=3.9952e-12 PD=1.012e-05 PS=1.992e-05 NRD=0.114537 NRS=0.193833 m=1 nf=2 $X=2590 $Y=4695 $D=8
XM5 a enb 12 vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=6280 $Y=5895 $D=8
X10 11 vdd ab vdd pmos_1p2_161 $T=3865 11540 1 0 $X=2435 $Y=9910
X11 12 11 en vdd pmos_1p2_161 $T=6435 11540 1 0 $X=5005 $Y=9910
.ENDS
***************************************
.SUBCKT M1_PSUB$$47335468
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT xpredec0_bot 1 2 3 8 9 10 11
** N=33 EP=7 IP=7 FDC=12
XM0 2 33 1 1 nfet_03v3 L=2.8e-07 W=3.285e-06 AD=3.0976e-12 AS=3.0976e-12 PD=1.496e-05 PS=1.496e-05 NRD=0.0625 NRS=0.0625 m=1 nf=1 $X=3755 $Y=35615 $D=2
XM1 3 2 1 1 nfet_03v3 L=2.8e-07 W=2.435e-06 AD=2.2968e-12 AS=2.2968e-12 PD=1.132e-05 PS=1.132e-05 NRD=0.0842912 NRS=0.0842912 m=1 nf=1 $X=6325 $Y=36010 $D=2
XM2 2 33 8 8 pfet_03v3 L=2.8e-07 W=8.255e-06 AD=7.7836e-12 AS=7.7836e-12 PD=3.626e-05 PS=3.626e-05 NRD=0.0248728 NRS=0.0248728 m=1 nf=1 $X=3755 $Y=16320 $D=8
XM3 3 2 8 8 pfet_03v3 L=2.8e-07 W=6.14e-06 AD=5.7904e-12 AS=5.7904e-12 PD=2.72e-05 PS=2.72e-05 NRD=0.0334347 NRS=0.0334347 m=1 nf=1 $X=6325 $Y=20855 $D=8
X4 1 33 9 8 11 10 alatch $T=350 -3160 0 0 $X=-100 $Y=-3165
.ENDS
***************************************
.SUBCKT xpredec0 vss vdd men clk A[1] A[0] x[3] x[2] x[1] x[0]
** N=99 EP=10 IP=158 FDC=56
XM0 x[3] 90 vss vss nfet_03v3 L=2.8e-07 W=8.47e-06 AD=4.7216e-12 AS=5.5388e-12 PD=2.024e-05 PS=2.514e-05 NRD=0.229075 NRS=0.268722 m=1 nf=4 $X=260 $Y=50820 $D=2
XM1 x[2] 92 vss vss nfet_03v3 L=2.8e-07 W=8.47e-06 AD=4.7216e-12 AS=4.7216e-12 PD=2.024e-05 PS=2.024e-05 NRD=0.229075 NRS=0.229075 m=1 nf=4 $X=4740 $Y=50820 $D=2
XM2 x[1] 94 vss vss nfet_03v3 L=2.8e-07 W=8.47e-06 AD=4.7216e-12 AS=4.7216e-12 PD=2.024e-05 PS=2.024e-05 NRD=0.229075 NRS=0.229075 m=1 nf=4 $X=9220 $Y=50820 $D=2
XM3 x[0] 96 vss vss nfet_03v3 L=2.8e-07 W=8.47e-06 AD=4.7216e-12 AS=5.5388e-12 PD=2.024e-05 PS=2.514e-05 NRD=0.229075 NRS=0.268722 m=1 nf=4 $X=13700 $Y=50820 $D=2
XM4 17 men vss vss nfet_03v3 L=2.8e-07 W=6.35e-07 AD=3.562e-13 AS=6.028e-13 PD=1.89e-06 PS=3.62e-06 NRD=0.189781 NRS=0.321168 m=1 nf=1 $X=21630 $Y=51200 $D=2
XM5 vss clk 17 vss nfet_03v3 L=2.8e-07 W=6.35e-07 AD=6.028e-13 AS=3.562e-13 PD=3.62e-06 PS=1.89e-06 NRD=0.321168 NRS=0.189781 m=1 nf=1 $X=22750 $Y=51200 $D=2
XM6 x[3] 90 vdd vdd pfet_03v3 L=2.8e-07 W=2.116e-05 AD=1.17936e-11 AS=1.38348e-11 PD=4.744e-05 PS=5.914e-05 NRD=0.0917108 NRS=0.107584 m=1 nf=4 $X=260 $Y=38080 $D=8
XM7 x[2] 92 vdd vdd pfet_03v3 L=2.8e-07 W=2.116e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.744e-05 PS=4.744e-05 NRD=0.0917108 NRS=0.0917108 m=1 nf=4 $X=4740 $Y=38080 $D=8
XM8 x[1] 94 vdd vdd pfet_03v3 L=2.8e-07 W=2.116e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.744e-05 PS=4.744e-05 NRD=0.0917108 NRS=0.0917108 m=1 nf=4 $X=9220 $Y=38080 $D=8
XM9 x[0] 96 vdd vdd pfet_03v3 L=2.8e-07 W=2.116e-05 AD=1.17936e-11 AS=1.38348e-11 PD=4.744e-05 PS=5.914e-05 NRD=0.0917108 NRS=0.107584 m=1 nf=4 $X=13700 $Y=38080 $D=8
XM10 98 men vdd vdd pfet_03v3 L=2.8e-07 W=7.95e-07 AD=4.39037e-13 AS=1.01447e-12 PD=2.22e-06 PS=4.6e-06 NRD=0.151026 NRS=0.348974 m=1 nf=1 $X=21630 $Y=47525 $D=8
XM11 17 clk 98 vdd pfet_03v3 L=2.8e-07 W=7.95e-07 AD=8.525e-15 AS=-8.525e-15 PD=1e-08 PS=-1e-08 NRD=0.00293255 NRS=-0.00293255 m=1 nf=1 $X=22745 $Y=47525 $D=8
XM12 99 clk 17 vdd pfet_03v3 L=2.8e-07 W=7.95e-07 AD=-8.525e-15 AS=8.525e-15 PD=-1e-08 PS=1e-08 NRD=-0.00293255 NRS=0.00293255 m=1 nf=1 $X=23870 $Y=47525 $D=8
XM13 vdd men 99 vdd pfet_03v3 L=2.8e-07 W=7.95e-07 AD=1.01447e-12 AS=4.39037e-13 PD=4.6e-06 PS=2.22e-06 NRD=0.348974 NRS=0.151026 m=1 nf=1 $X=24985 $Y=47525 $D=8
XM14 18 17 vdd vdd pfet_03v3 L=2.8e-07 W=1.06e-06 AD=5.928e-13 AS=1.0032e-12 PD=3.32e-06 PS=6.32e-06 NRD=0.45614 NRS=0.77193 m=1 nf=2 $X=29010 $Y=47595 $D=8
X17 18 vss 17 vss nmos_1p2$$46563372 $T=29755 51180 0 0 $X=28610 $Y=50495
X18 90 vss vdd 30 31 xpredec0_xa $T=-2205 170 0 0 $X=-1440 $Y=-5
X19 92 vss vdd 30 32 xpredec0_xa $T=11165 170 1 180 $X=3000 $Y=-5
X20 94 vss vdd 33 31 xpredec0_xa $T=6755 170 0 0 $X=7520 $Y=-5
X21 96 vss vdd 33 32 xpredec0_xa $T=20125 170 1 180 $X=11960 $Y=-5
X22 vss 30 33 vdd A[1] 17 18 xpredec0_bot $T=18665 3160 0 0 $X=18135 $Y=-5
X23 vss 31 32 vdd A[0] 17 18 xpredec0_bot $T=27120 3160 0 0 $X=26590 $Y=-5
.ENDS
***************************************
.SUBCKT M1_PACTIVE_I02
** N=38 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pfet_03v3_I01
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_03v3_I04
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ypredec1_ys
** N=8 EP=0 IP=36 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_32 1 2 4 5 7 8
** N=8 EP=6 IP=10 FDC=4
*.SEEDPROM
XM0 1 7 4 1 nfet_03v3 L=2.8e-07 W=1.271e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=3510 $Y=1700 $D=2
XM1 8 5 1 1 nfet_03v3 L=2.8e-07 W=4.235e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=6870 $Y=1700 $D=2
XM2 2 7 4 2 pfet_03v3 L=2.8e-07 W=2.8e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=3510 $Y=14855 $D=8
XM3 8 5 2 2 pfet_03v3 L=2.8e-07 W=9.33e-06 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=6870 $Y=14855 $D=8
.ENDS
***************************************
.SUBCKT ICV_33 1 2 4 5 6 7 8 9 11 13
** N=14 EP=10 IP=16 FDC=12
*.SEEDPROM
XM0 1 14 6 1 nfet_03v3 L=2.8e-07 W=1.271e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=9110 $Y=1700 $D=2
XM1 12 7 1 1 nfet_03v3 L=2.8e-07 W=4.235e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=12470 $Y=1700 $D=2
XM2 2 14 6 2 pfet_03v3 L=2.8e-07 W=2.8e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=9110 $Y=14855 $D=8
XM3 12 7 2 2 pfet_03v3 L=2.8e-07 W=9.33e-06 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=12470 $Y=14855 $D=8
X4 1 2 4 5 11 14 ICV_32 $T=0 0 0 0 $X=-5 $Y=-5
X5 1 2 8 9 12 13 ICV_32 $T=11200 0 0 0 $X=11195 $Y=-5
.ENDS
***************************************
.SUBCKT nmos_1p2$$47514668
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ypredec1_bot 1 2 3 10 11 12 13
** N=34 EP=7 IP=20 FDC=12
XM0 2 30 1 1 nfet_03v3 L=2.8e-07 W=2.115e-06 AD=1.9976e-12 AS=1.9976e-12 PD=9.96e-06 PS=9.96e-06 NRD=0.0969163 NRS=0.0969163 m=1 nf=1 $X=3755 $Y=33350 $D=2
XM1 3 2 1 1 nfet_03v3 L=2.8e-07 W=2.115e-06 AD=1.9976e-12 AS=1.9976e-12 PD=9.96e-06 PS=9.96e-06 NRD=0.0969163 NRS=0.0969163 m=1 nf=1 $X=6325 $Y=33350 $D=2
X2 10 2 30 pmos_1p2$$46887980 $T=3910 18340 0 0 $X=2480 $Y=17630
X3 10 3 2 pmos_1p2$$46887980 $T=6480 18340 0 0 $X=5050 $Y=17630
X4 1 30 11 10 13 12 alatch $T=350 -3160 0 0 $X=-100 $Y=-3165
.ENDS
***************************************
.SUBCKT pmos_1p2$$47821868
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$47820844
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ypredec1_xa
** N=29 EP=0 IP=36 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_34 1 2 5 8 9 10 11 12
** N=22 EP=8 IP=36 FDC=16
XM0 20 10 13 1 nfet_03v3 L=2.8e-07 W=3.175e-06 AD=1.73655e-12 AS=4.05195e-12 PD=7.32e-06 PS=1.481e-05 NRD=0.0374449 NRS=0.0873715 m=1 nf=1 $X=-2370 $Y=-33035 $D=2
XM1 19 9 20 1 nfet_03v3 L=2.8e-07 W=3.175e-06 AD=3.405e-14 AS=-3.405e-14 PD=1e-08 PS=-1e-08 NRD=0.000734214 NRS=-0.000734214 m=1 nf=1 $X=-1260 $Y=-33035 $D=2
XM2 1 2 19 1 nfet_03v3 L=2.8e-07 W=3.175e-06 AD=3.405e-14 AS=-3.405e-14 PD=1e-08 PS=-1e-08 NRD=0.000734214 NRS=-0.000734214 m=1 nf=1 $X=-140 $Y=-33035 $D=2
XM3 1 13 11 1 nfet_03v3 L=2.8e-07 W=3.175e-06 AD=1.7706e-12 AS=2.1792e-12 PD=8.37e-06 PS=1.1e-05 NRD=0.343612 NRS=0.422907 m=1 nf=3 $X=-2375 $Y=-2950 $D=2
XM4 21 5 1 1 nfet_03v3 L=2.8e-07 W=3.175e-06 AD=-3.405e-14 AS=3.405e-14 PD=-1e-08 PS=1e-08 NRD=-0.000734214 NRS=0.000734214 m=1 nf=1 $X=990 $Y=-33035 $D=2
XM5 22 9 21 1 nfet_03v3 L=2.8e-07 W=3.175e-06 AD=-3.405e-14 AS=3.405e-14 PD=-1e-08 PS=1e-08 NRD=-0.000734214 NRS=0.000734214 m=1 nf=1 $X=2110 $Y=-33035 $D=2
XM6 16 10 22 1 nfet_03v3 L=2.8e-07 W=3.175e-06 AD=4.05195e-12 AS=1.73655e-12 PD=1.481e-05 PS=7.32e-06 NRD=0.0873715 NRS=0.0374449 m=1 nf=1 $X=3220 $Y=-33035 $D=2
XM7 12 16 1 1 nfet_03v3 L=2.8e-07 W=3.175e-06 AD=2.1792e-12 AS=1.7706e-12 PD=1.1e-05 PS=8.37e-06 NRD=0.422907 NRS=0.343612 m=1 nf=3 $X=985 $Y=-2950 $D=2
XM8 8 10 13 8 pfet_03v3 L=2.8e-07 W=2.645e-06 AD=1.4742e-12 AS=2.4948e-12 PD=6.19e-06 PS=1.222e-05 NRD=0.0458554 NRS=0.0776014 m=1 nf=1 $X=-2375 $Y=-19360 $D=8
XM9 13 9 8 8 pfet_03v3 L=2.8e-07 W=2.645e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=-1255 $Y=-19360 $D=8
XM10 8 2 13 8 pfet_03v3 L=2.8e-07 W=2.645e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=-135 $Y=-19360 $D=8
XM11 8 13 11 8 pfet_03v3 L=2.8e-07 W=8.075e-06 AD=4.5006e-12 AS=5.5392e-12 PD=1.887e-05 PS=2.5e-05 NRD=0.135182 NRS=0.166378 m=1 nf=3 $X=-2375 $Y=-10125 $D=8
XM12 16 5 8 8 pfet_03v3 L=2.8e-07 W=2.645e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=985 $Y=-19360 $D=8
XM13 8 9 16 8 pfet_03v3 L=2.8e-07 W=2.645e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=2105 $Y=-19360 $D=8
XM14 16 10 8 8 pfet_03v3 L=2.8e-07 W=2.645e-06 AD=2.4948e-12 AS=1.4742e-12 PD=1.222e-05 PS=6.19e-06 NRD=0.0776014 NRS=0.0458554 m=1 nf=1 $X=3225 $Y=-19360 $D=8
XM15 12 16 8 8 pfet_03v3 L=2.8e-07 W=8.075e-06 AD=5.5392e-12 AS=4.5006e-12 PD=2.5e-05 PS=1.887e-05 NRD=0.166378 NRS=0.135182 m=1 nf=3 $X=985 $Y=-10125 $D=8
.ENDS
***************************************
.SUBCKT pmos_1p2$$47109164 1 2 3
** N=4 EP=3 IP=0 FDC=1
XM0 2 3 1 1 pfet_03v3 L=2.8e-07 W=1.595e-06 AD=8.892e-13 AS=1.5048e-12 PD=4.46e-06 PS=8.6e-06 NRD=0.304094 NRS=0.51462 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nmos_1p2$$47342636
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_03v3_I18
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ypredec1 1 2 men clk ly[6] ly[7] ly[0] ly[1] ly[2] ly[3] ly[4] ly[5] ry[0] ry[1] ry[2] ry[3] ry[4] ry[5] ry[6] ry[7]
+ A[2] A[1] A[0]
** N=374 EP=23 IP=151 FDC=172
XM0 367 358 1 1 nfet_03v3 L=2.8e-07 W=4.235e-06 AD=3.9952e-12 AS=3.9952e-12 PD=1.904e-05 PS=1.904e-05 NRD=0.0484581 NRS=0.0484581 m=1 nf=1 $X=2545 $Y=46970 $D=2
XM1 1 371 ly[3] 1 nfet_03v3 L=2.8e-07 W=1.271e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=21585 $Y=46970 $D=2
XM2 368 361 1 1 nfet_03v3 L=2.8e-07 W=4.235e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=24945 $Y=46970 $D=2
XM3 188 189 1 1 nfet_03v3 L=2.8e-07 W=6.3e-07 AD=5.984e-13 AS=5.984e-13 PD=3.6e-06 PS=3.6e-06 NRD=0.323529 NRS=0.323529 m=1 nf=1 $X=31760 $Y=4985 $D=2
XM4 189 clk 1 1 nfet_03v3 L=2.8e-07 W=8.9e-07 AD=4.966e-13 AS=8.404e-13 PD=2.43e-06 PS=4.7e-06 NRD=0.136126 NRS=0.230366 m=1 nf=1 $X=38610 $Y=5010 $D=2
XM5 1 men 189 1 nfet_03v3 L=2.8e-07 W=8.9e-07 AD=8.404e-13 AS=4.966e-13 PD=4.7e-06 PS=2.43e-06 NRD=0.230366 NRS=0.136126 m=1 nf=1 $X=39730 $Y=5010 $D=2
XM6 1 372 ly[7] 1 nfet_03v3 L=2.8e-07 W=1.271e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=43985 $Y=46970 $D=2
XM7 369 358 1 1 nfet_03v3 L=2.8e-07 W=4.235e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=47345 $Y=46970 $D=2
XM8 1 373 ry[3] 1 nfet_03v3 L=2.8e-07 W=1.271e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=66385 $Y=46970 $D=2
XM9 370 361 1 1 nfet_03v3 L=2.8e-07 W=4.235e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=69745 $Y=46970 $D=2
XM10 1 374 ry[7] 1 nfet_03v3 L=2.8e-07 W=1.271e-05 AD=8.7168e-12 AS=8.7168e-12 PD=3.824e-05 PS=3.824e-05 NRD=0.105727 NRS=0.105727 m=1 nf=3 $X=88785 $Y=46970 $D=2
XM11 367 358 2 2 pfet_03v3 L=2.8e-07 W=9.33e-06 AD=8.8e-12 AS=8.8e-12 PD=4.088e-05 PS=4.088e-05 NRD=0.022 NRS=0.022 m=1 nf=1 $X=2545 $Y=60125 $D=8
XM12 2 371 ly[3] 2 pfet_03v3 L=2.8e-07 W=2.8e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=21585 $Y=60125 $D=8
XM13 368 361 2 2 pfet_03v3 L=2.8e-07 W=9.33e-06 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=24945 $Y=60125 $D=8
XM14 365 men 2 2 pfet_03v3 L=2.8e-07 W=1.06e-06 AD=5.915e-13 AS=1.35362e-12 PD=2.795e-06 PS=5.74e-06 NRD=0.114286 NRS=0.261538 m=1 nf=1 $X=36375 $Y=1335 $D=8
XM15 189 clk 365 2 pfet_03v3 L=2.8e-07 W=1.06e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=37495 $Y=1335 $D=8
XM16 366 clk 189 2 pfet_03v3 L=2.8e-07 W=1.06e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=38615 $Y=1335 $D=8
XM17 2 men 366 2 pfet_03v3 L=2.8e-07 W=1.06e-06 AD=1.34225e-12 AS=5.915e-13 PD=5.73e-06 PS=2.795e-06 NRD=0.259341 NRS=0.114286 m=1 nf=1 $X=39735 $Y=1335 $D=8
XM18 2 372 ly[7] 2 pfet_03v3 L=2.8e-07 W=2.8e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=43985 $Y=60125 $D=8
XM19 369 358 2 2 pfet_03v3 L=2.8e-07 W=9.33e-06 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=47345 $Y=60125 $D=8
XM20 2 373 ry[3] 2 pfet_03v3 L=2.8e-07 W=2.8e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=66385 $Y=60125 $D=8
XM21 370 361 2 2 pfet_03v3 L=2.8e-07 W=9.33e-06 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=69745 $Y=60125 $D=8
XM22 2 374 ry[7] 2 pfet_03v3 L=2.8e-07 W=2.8e-05 AD=1.92e-11 AS=1.92e-11 PD=8.192e-05 PS=8.192e-05 NRD=0.048 NRS=0.048 m=1 nf=3 $X=88785 $Y=60125 $D=8
X23 1 2 ly[0] 357 ly[1] 359 ly[2] 360 367 371 ICV_33 $T=1275 45270 0 0 $X=1270 $Y=45265
X24 1 2 ly[4] 362 ly[5] 363 ly[6] 364 368 372 ICV_33 $T=23675 45270 0 0 $X=23670 $Y=45265
X25 1 2 ry[0] 357 ry[1] 359 ry[2] 360 369 373 ICV_33 $T=46075 45270 0 0 $X=46070 $Y=45265
X26 1 2 ry[4] 362 ry[5] 363 ry[6] 364 370 374 ICV_33 $T=68475 45270 0 0 $X=68470 $Y=45265
X27 1 190 191 2 A[2] 189 188 ypredec1_bot $T=1920 5135 0 0 $X=1820 $Y=1970
X28 1 192 193 2 A[1] 189 188 ypredec1_bot $T=10375 5135 0 0 $X=10275 $Y=1970
X29 1 194 195 2 A[0] 189 188 ypredec1_bot $T=18830 5135 0 0 $X=18730 $Y=1970
X30 1 195 194 2 192 190 363 364 ICV_34 $T=33645 42985 1 180 $X=28115 $Y=7365
X31 1 195 194 2 193 190 361 362 ICV_34 $T=41810 42985 1 180 $X=36280 $Y=7365
X32 1 195 194 2 192 191 359 360 ICV_34 $T=49980 42985 1 180 $X=44450 $Y=7365
X33 1 195 194 2 193 191 358 357 ICV_34 $T=58150 42985 1 180 $X=52620 $Y=7365
X34 2 188 189 pmos_1p2$$47109164 $T=32795 1405 1 180 $X=28795 $Y=720
.ENDS
***************************************
.SUBCKT M1_NWELL_01
** N=49 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nfet_03v3_I20 1 2 3
** N=3 EP=3 IP=0 FDC=1
XM0 2 3 1 2 nfet_03v3 L=2.8e-07 W=4.715e-06 AD=4.4484e-12 AS=4.4484e-12 PD=2.11e-05 PS=2.11e-05 NRD=0.0435213 NRS=0.0435213 m=1 nf=1 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT M1_PACTIVE$10
** N=13 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pmos_1p2_02_R90 1 2 3
** N=3 EP=3 IP=0 FDC=1
XM0 2 3 1 1 pfet_03v3 L=2.8e-07 W=1.178e-05 AD=6.5676e-12 AS=1.11144e-11 PD=2.63e-05 PS=5.228e-05 NRD=0.0411718 NRS=0.0696754 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pfet_03v3_I14 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
XM0 2 3 1 4 pfet_03v3 L=2.8e-07 W=3.075e-06 AD=2.8996e-12 AS=2.8996e-12 PD=1.406e-05 PS=1.406e-05 NRD=0.0667678 NRS=0.0667678 m=1 nf=1 $X=0 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nfet_03v3_I11 1 2 3
** N=3 EP=3 IP=0 FDC=1
XM0 2 3 1 2 nfet_03v3 L=2.8e-07 W=1.23e-06 AD=1.1616e-12 AS=1.1616e-12 PD=6.16e-06 PS=6.16e-06 NRD=0.166667 NRS=0.166667 m=1 nf=1 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pfet_03v3_I17 1 2 3
** N=3 EP=3 IP=0 FDC=1
XM0 2 3 1 1 pfet_03v3 L=2.8e-07 W=2.203e-05 AD=1.2272e-11 AS=1.39712e-11 PD=5.24e-05 PS=6.256e-05 NRD=0.550847 NRS=0.627119 m=1 nf=10 $X=0 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nfet_03v3_I06 1 2 3
** N=3 EP=3 IP=0 FDC=1
XM0 2 3 1 1 nfet_03v3 L=2.8e-07 W=8.96e-06 AD=4.992e-12 AS=5.6832e-12 PD=2.44e-05 PS=2.896e-05 NRD=1.35417 NRS=1.54167 m=1 nf=10 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT M1_PACTIVE_I01
** N=7 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT wen_v2 vss vdd wen clk IGWEN GWE
** N=50 EP=6 IP=93 FDC=30
XM0 vss wen 28 vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=2545 $Y=1065 $D=2
XM1 11 wen vss vss nfet_03v3 L=2.8e-07 W=2.8e-06 AD=1.92e-12 AS=1.92e-12 PD=9.92e-06 PS=9.92e-06 NRD=0.48 NRS=0.48 m=1 nf=3 $X=1260 $Y=16070 $D=2
XM2 29 clk vss vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=3665 $Y=1065 $D=2
XM3 30 29 vss vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=5905 $Y=1475 $D=2
XM4 33 29 28 vss nfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=8440 $Y=545 $D=2
XM5 34 30 33 vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=10750 $Y=1860 $D=2
XM6 vss 35 34 vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=11870 $Y=1860 $D=2
XM7 vss 33 35 vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=14110 $Y=1860 $D=2
XM8 15 35 vss vss nfet_03v3 L=2.8e-07 W=1.12e-06 AD=6.24e-13 AS=1.056e-12 PD=3.44e-06 PS=6.56e-06 NRD=0.433333 NRS=0.733333 m=1 nf=2 $X=16465 $Y=1620 $D=2
XM9 15 30 31 vss nfet_03v3 L=2.8e-07 W=2.115e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=19750 $Y=545 $D=2
XM10 32 29 31 vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=23090 $Y=1240 $D=2
XM11 vss 19 32 vss nfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=24210 $Y=1240 $D=2
XM12 19 31 vss vss nfet_03v3 L=2.8e-07 W=2.905e-06 AD=1.78e-12 AS=1.78e-12 PD=1.112e-05 PS=1.112e-05 NRD=2.24719 NRS=2.24719 m=1 nf=7 $X=26535 $Y=1905 $D=2
XM13 vdd wen 28 vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=2545 $Y=4215 $D=8
XM14 29 clk vdd vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=3665 $Y=4215 $D=8
XM15 30 29 vdd vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=5905 $Y=4215 $D=8
XM16 11 wen vdd vdd pfet_03v3 L=2.8e-07 W=6.94e-06 AD=3.8688e-12 AS=4.7616e-12 PD=1.8e-05 PS=2.368e-05 NRD=0.629032 NRS=0.774194 m=1 nf=6 $X=1260 $Y=9420 $D=8
XM17 33 30 28 vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=1.17422e-12 AS=9.988e-13 PD=4.793e-06 PS=5.42e-06 NRD=0.227875 NRS=0.193833 m=1 nf=1 $X=8440 $Y=4215 $D=8
XM18 34 29 33 vdd pfet_03v3 L=2.8e-07 W=4.45e-07 AD=-6.91897e-13 AS=-6.43897e-13 PD=-2.79573e-06 PS=-2.69573e-06 NRD=-0.750757 NRS=-0.698673 m=1 nf=1 $X=10180 $Y=4215 $D=8
XM19 vdd 35 34 vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=1.14048e-12 PD=5.42e-06 PS=4.72272e-06 NRD=0.193833 NRS=0.221328 m=1 nf=1 $X=11870 $Y=4215 $D=8
XM20 vdd 33 35 vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=14110 $Y=4215 $D=8
XM21 15 35 vdd vdd pfet_03v3 L=2.8e-07 W=2.65e-06 AD=1.4768e-12 AS=2.4992e-12 PD=6.72e-06 PS=1.312e-05 NRD=0.183099 NRS=0.309859 m=1 nf=2 $X=16465 $Y=4215 $D=8
XM22 15 29 31 vdd pfet_03v3 L=2.8e-07 W=2.115e-06 AD=1.1804e-12 AS=2.13253e-12 PD=5.58e-06 PS=1.01287e-05 NRD=0.229075 NRS=0.413851 m=1 nf=2 $X=19750 $Y=4215 $D=8
XM23 32 30 31 vdd pfet_03v3 L=2.8e-07 W=4.45e-07 AD=-6.59976e-13 AS=-6.40776e-13 PD=-2.72923e-06 PS=-2.68923e-06 NRD=-0.71612 NRS=-0.695287 m=1 nf=1 $X=22550 $Y=5525 $D=8
XM24 vdd 19 32 vdd pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=1.12024e-12 PD=5.42e-06 PS=4.68056e-06 NRD=0.193833 NRS=0.2174 m=1 nf=1 $X=24210 $Y=4215 $D=8
XM25 19 31 vdd vdd pfet_03v3 L=2.8e-07 W=7.185e-06 AD=4.4e-12 AS=4.4e-12 PD=2.16e-05 PS=2.16e-05 NRD=0.909091 NRS=0.909091 m=1 nf=7 $X=26535 $Y=4215 $D=8
X46 vdd IGWEN 11 pfet_03v3_I17 $T=10115 9420 0 0 $X=9075 $Y=8800
X47 vdd GWE 19 pfet_03v3_I17 $T=23345 9420 0 0 $X=22305 $Y=8800
X48 vss IGWEN 11 nfet_03v3_I06 $T=10115 16070 0 0 $X=9435 $Y=15450
X49 vss GWE 19 nfet_03v3_I06 $T=23345 16070 0 0 $X=22665 $Y=15450
.ENDS
***************************************
.SUBCKT pmos_1p2$$47512620
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT xpredec1_xa
** N=29 EP=0 IP=36 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$47337516 1 2 3
** N=3 EP=3 IP=0 FDC=1
XM0 2 3 1 1 pfet_03v3 L=2.8e-07 W=7.62e-06 AD=7.1852e-12 AS=7.1852e-12 PD=3.354e-05 PS=3.354e-05 NRD=0.0269443 NRS=0.0269443 m=1 nf=1 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nmos_1p2$$47336492 1 2 3
** N=3 EP=3 IP=0 FDC=1
XM0 2 3 1 1 nfet_03v3 L=2.8e-07 W=3.07e-06 AD=2.8952e-12 AS=2.8952e-12 PD=1.404e-05 PS=1.404e-05 NRD=0.0668693 NRS=0.0668693 m=1 nf=1 $X=-155 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT xpredec1_bot 1 2 3 10 11 12 13
** N=32 EP=7 IP=19 FDC=12
X0 1 32 11 10 13 12 alatch $T=350 -3160 0 0 $X=-100 $Y=-3165
X2 10 2 32 pmos_1p2$$47337516 $T=3910 18340 0 0 $X=2480 $Y=17635
X3 10 3 2 pmos_1p2$$47337516 $T=6480 18340 0 0 $X=5050 $Y=17635
X4 1 2 32 nmos_1p2$$47336492 $T=3910 36070 0 0 $X=2765 $Y=35385
X5 1 3 2 nmos_1p2$$47336492 $T=6480 36070 0 0 $X=5335 $Y=35385
.ENDS
***************************************
.SUBCKT xpredec1 vss men vdd clk A[2] A[1] A[0] x[7] x[6] x[5] x[4] x[3] x[2] x[1] x[0]
** N=91 EP=15 IP=199 FDC=108
XM0 77 18 51 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=3.2435e-12 AS=7.36025e-12 PD=1.2995e-05 PS=2.613e-05 NRD=0.0208417 NRS=0.0472946 m=1 nf=1 $X=1700 $Y=2310 $D=2
XM1 76 19 77 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=2820 $Y=2310 $D=2
XM2 vss 20 76 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=3940 $Y=2310 $D=2
XM3 vss 51 x[7] vss nfet_03v3 L=2.8e-07 W=6.355e-06 AD=3.5412e-12 AS=4.3584e-12 PD=1.518e-05 PS=2.008e-05 NRD=0.171806 NRS=0.211454 m=1 nf=3 $X=1700 $Y=48000 $D=2
XM4 78 21 vss vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=5060 $Y=2310 $D=2
XM5 79 19 78 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=6180 $Y=2310 $D=2
XM6 54 18 79 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=7.36025e-12 AS=3.2435e-12 PD=2.613e-05 PS=1.2995e-05 NRD=0.0472946 NRS=0.0208417 m=1 nf=1 $X=7300 $Y=2310 $D=2
XM7 x[6] 54 vss vss nfet_03v3 L=2.8e-07 W=6.355e-06 AD=4.3584e-12 AS=3.5412e-12 PD=2.008e-05 PS=1.518e-05 NRD=0.211454 NRS=0.171806 m=1 nf=3 $X=5060 $Y=48000 $D=2
XM8 81 18 57 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=3.2435e-12 AS=7.36025e-12 PD=1.2995e-05 PS=2.613e-05 NRD=0.0208417 NRS=0.0472946 m=1 nf=1 $X=9870 $Y=2310 $D=2
XM9 80 22 81 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=10990 $Y=2310 $D=2
XM10 vss 20 80 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=12110 $Y=2310 $D=2
XM11 vss 57 x[5] vss nfet_03v3 L=2.8e-07 W=6.355e-06 AD=3.5412e-12 AS=4.3584e-12 PD=1.518e-05 PS=2.008e-05 NRD=0.171806 NRS=0.211454 m=1 nf=3 $X=9870 $Y=48000 $D=2
XM12 82 21 vss vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=13230 $Y=2310 $D=2
XM13 83 22 82 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=14350 $Y=2310 $D=2
XM14 60 18 83 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=7.36025e-12 AS=3.2435e-12 PD=2.613e-05 PS=1.2995e-05 NRD=0.0472946 NRS=0.0208417 m=1 nf=1 $X=15470 $Y=2310 $D=2
XM15 x[4] 60 vss vss nfet_03v3 L=2.8e-07 W=6.355e-06 AD=4.3584e-12 AS=3.5412e-12 PD=2.008e-05 PS=1.518e-05 NRD=0.211454 NRS=0.171806 m=1 nf=3 $X=13230 $Y=48000 $D=2
XM16 85 23 63 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=3.2435e-12 AS=7.36025e-12 PD=1.2995e-05 PS=2.613e-05 NRD=0.0208417 NRS=0.0472946 m=1 nf=1 $X=18035 $Y=2310 $D=2
XM17 84 19 85 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=19155 $Y=2310 $D=2
XM18 vss 20 84 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=20275 $Y=2310 $D=2
XM19 vss 63 x[3] vss nfet_03v3 L=2.8e-07 W=6.355e-06 AD=3.5412e-12 AS=4.3584e-12 PD=1.518e-05 PS=2.008e-05 NRD=0.171806 NRS=0.211454 m=1 nf=3 $X=18035 $Y=48000 $D=2
XM20 86 21 vss vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=21395 $Y=2310 $D=2
XM21 87 19 86 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=22515 $Y=2310 $D=2
XM22 66 23 87 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=7.36025e-12 AS=3.2435e-12 PD=2.613e-05 PS=1.2995e-05 NRD=0.0472946 NRS=0.0208417 m=1 nf=1 $X=23635 $Y=2310 $D=2
XM23 x[2] 66 vss vss nfet_03v3 L=2.8e-07 W=6.355e-06 AD=4.3584e-12 AS=3.5412e-12 PD=2.008e-05 PS=1.518e-05 NRD=0.211454 NRS=0.171806 m=1 nf=3 $X=21395 $Y=48000 $D=2
XM24 89 23 69 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=3.2435e-12 AS=7.36025e-12 PD=1.2995e-05 PS=2.613e-05 NRD=0.0208417 NRS=0.0472946 m=1 nf=1 $X=26205 $Y=2310 $D=2
XM25 88 22 89 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=27325 $Y=2310 $D=2
XM26 vss 20 88 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=28445 $Y=2310 $D=2
XM27 vss 69 x[1] vss nfet_03v3 L=2.8e-07 W=6.355e-06 AD=3.5412e-12 AS=4.3584e-12 PD=1.518e-05 PS=2.008e-05 NRD=0.171806 NRS=0.211454 m=1 nf=3 $X=26205 $Y=48000 $D=2
XM28 90 21 vss vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=29565 $Y=2310 $D=2
XM29 91 22 90 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=30685 $Y=2310 $D=2
XM30 72 23 91 vss nfet_03v3 L=2.8e-07 W=5.82e-06 AD=7.36025e-12 AS=3.2435e-12 PD=2.613e-05 PS=1.2995e-05 NRD=0.0472946 NRS=0.0208417 m=1 nf=1 $X=31805 $Y=2310 $D=2
XM31 x[0] 72 vss vss nfet_03v3 L=2.8e-07 W=6.355e-06 AD=4.3584e-12 AS=3.5412e-12 PD=2.008e-05 PS=1.518e-05 NRD=0.211454 NRS=0.171806 m=1 nf=3 $X=29565 $Y=48000 $D=2
XM32 17 men vss vss nfet_03v3 L=2.8e-07 W=8.9e-07 AD=4.966e-13 AS=8.404e-13 PD=2.43e-06 PS=4.7e-06 NRD=0.136126 NRS=0.230366 m=1 nf=1 $X=37165 $Y=51200 $D=2
XM33 vss clk 17 vss nfet_03v3 L=2.8e-07 W=8.9e-07 AD=8.404e-13 AS=4.966e-13 PD=4.7e-06 PS=2.43e-06 NRD=0.230366 NRS=0.136126 m=1 nf=1 $X=38285 $Y=51200 $D=2
XM34 vss 17 16 vss nfet_03v3 L=2.8e-07 W=6.3e-07 AD=5.984e-13 AS=5.984e-13 PD=3.6e-06 PS=3.6e-06 NRD=0.323529 NRS=0.323529 m=1 nf=1 $X=45140 $Y=51180 $D=2
XM35 vdd 18 51 vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=2.7118e-12 AS=4.5892e-12 PD=1.095e-05 PS=2.174e-05 NRD=0.0249281 NRS=0.042186 m=1 nf=1 $X=1700 $Y=21650 $D=8
XM36 51 19 vdd vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=2820 $Y=21650 $D=8
XM37 vdd 20 51 vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=3940 $Y=21650 $D=8
XM38 vdd 51 x[7] vdd pfet_03v3 L=2.8e-07 W=1.587e-05 AD=8.8452e-12 AS=1.08864e-11 PD=3.558e-05 PS=4.728e-05 NRD=0.0687831 NRS=0.0846561 m=1 nf=3 $X=1700 $Y=35260 $D=8
XM39 54 21 vdd vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=5060 $Y=21650 $D=8
XM40 vdd 19 54 vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=6180 $Y=21650 $D=8
XM41 54 18 vdd vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=4.5892e-12 AS=2.7118e-12 PD=2.174e-05 PS=1.095e-05 NRD=0.042186 NRS=0.0249281 m=1 nf=1 $X=7300 $Y=21650 $D=8
XM42 x[6] 54 vdd vdd pfet_03v3 L=2.8e-07 W=1.587e-05 AD=1.08864e-11 AS=8.8452e-12 PD=4.728e-05 PS=3.558e-05 NRD=0.0846561 NRS=0.0687831 m=1 nf=3 $X=5060 $Y=35260 $D=8
XM43 vdd 18 57 vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=2.7118e-12 AS=4.5892e-12 PD=1.095e-05 PS=2.174e-05 NRD=0.0249281 NRS=0.042186 m=1 nf=1 $X=9870 $Y=21650 $D=8
XM44 57 22 vdd vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=10990 $Y=21650 $D=8
XM45 vdd 20 57 vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=12110 $Y=21650 $D=8
XM46 vdd 57 x[5] vdd pfet_03v3 L=2.8e-07 W=1.587e-05 AD=8.8452e-12 AS=1.08864e-11 PD=3.558e-05 PS=4.728e-05 NRD=0.0687831 NRS=0.0846561 m=1 nf=3 $X=9870 $Y=35260 $D=8
XM47 60 21 vdd vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=13230 $Y=21650 $D=8
XM48 vdd 22 60 vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=14350 $Y=21650 $D=8
XM49 60 18 vdd vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=4.5892e-12 AS=2.7118e-12 PD=2.174e-05 PS=1.095e-05 NRD=0.042186 NRS=0.0249281 m=1 nf=1 $X=15470 $Y=21650 $D=8
XM50 x[4] 60 vdd vdd pfet_03v3 L=2.8e-07 W=1.587e-05 AD=1.08864e-11 AS=8.8452e-12 PD=4.728e-05 PS=3.558e-05 NRD=0.0846561 NRS=0.0687831 m=1 nf=3 $X=13230 $Y=35260 $D=8
XM51 vdd 23 63 vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=2.7118e-12 AS=4.5892e-12 PD=1.095e-05 PS=2.174e-05 NRD=0.0249281 NRS=0.042186 m=1 nf=1 $X=18035 $Y=21650 $D=8
XM52 63 19 vdd vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=19155 $Y=21650 $D=8
XM53 vdd 20 63 vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=20275 $Y=21650 $D=8
XM54 vdd 63 x[3] vdd pfet_03v3 L=2.8e-07 W=1.587e-05 AD=8.8452e-12 AS=1.08864e-11 PD=3.558e-05 PS=4.728e-05 NRD=0.0687831 NRS=0.0846561 m=1 nf=3 $X=18035 $Y=35260 $D=8
XM55 66 21 vdd vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=21395 $Y=21650 $D=8
XM56 vdd 19 66 vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=22515 $Y=21650 $D=8
XM57 66 23 vdd vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=4.5892e-12 AS=2.7118e-12 PD=2.174e-05 PS=1.095e-05 NRD=0.042186 NRS=0.0249281 m=1 nf=1 $X=23635 $Y=21650 $D=8
XM58 x[2] 66 vdd vdd pfet_03v3 L=2.8e-07 W=1.587e-05 AD=1.08864e-11 AS=8.8452e-12 PD=4.728e-05 PS=3.558e-05 NRD=0.0846561 NRS=0.0687831 m=1 nf=3 $X=21395 $Y=35260 $D=8
XM59 vdd 23 69 vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=2.7118e-12 AS=4.5892e-12 PD=1.095e-05 PS=2.174e-05 NRD=0.0249281 NRS=0.042186 m=1 nf=1 $X=26205 $Y=21650 $D=8
XM60 69 22 vdd vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=27325 $Y=21650 $D=8
XM61 vdd 20 69 vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=28445 $Y=21650 $D=8
XM62 vdd 69 x[1] vdd pfet_03v3 L=2.8e-07 W=1.587e-05 AD=8.8452e-12 AS=1.08864e-11 PD=3.558e-05 PS=4.728e-05 NRD=0.0687831 NRS=0.0846561 m=1 nf=3 $X=26205 $Y=35260 $D=8
XM63 72 21 vdd vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=29565 $Y=21650 $D=8
XM64 vdd 22 72 vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=30685 $Y=21650 $D=8
XM65 72 23 vdd vdd pfet_03v3 L=2.8e-07 W=4.865e-06 AD=4.5892e-12 AS=2.7118e-12 PD=2.174e-05 PS=1.095e-05 NRD=0.042186 NRS=0.0249281 m=1 nf=1 $X=31805 $Y=21650 $D=8
XM66 x[0] 72 vdd vdd pfet_03v3 L=2.8e-07 W=1.587e-05 AD=1.08864e-11 AS=8.8452e-12 PD=4.728e-05 PS=3.558e-05 NRD=0.0846561 NRS=0.0687831 m=1 nf=3 $X=29565 $Y=35260 $D=8
XM67 74 men vdd vdd pfet_03v3 L=2.8e-07 W=1.06e-06 AD=5.915e-13 AS=1.35362e-12 PD=2.795e-06 PS=5.74e-06 NRD=0.114286 NRS=0.261538 m=1 nf=1 $X=37165 $Y=47525 $D=8
XM68 17 clk 74 vdd pfet_03v3 L=2.8e-07 W=1.06e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=38285 $Y=47525 $D=8
XM69 75 clk 17 vdd pfet_03v3 L=2.8e-07 W=1.06e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=39405 $Y=47525 $D=8
XM70 vdd men 75 vdd pfet_03v3 L=2.8e-07 W=1.06e-06 AD=1.35362e-12 AS=5.915e-13 PD=5.74e-06 PS=2.795e-06 NRD=0.261538 NRS=0.114286 m=1 nf=1 $X=40525 $Y=47525 $D=8
X71 vdd 16 17 pmos_1p2$$47109164 $T=44700 47595 0 0 $X=42105 $Y=46910
X83 vss 18 23 vdd A[2] 17 16 xpredec1_bot $T=34205 3160 0 0 $X=33675 $Y=-5
X84 vss 19 22 vdd A[1] 17 16 xpredec1_bot $T=42655 3160 0 0 $X=42125 $Y=-5
X85 vss 20 21 vdd A[0] 17 16 xpredec1_bot $T=51110 3160 0 0 $X=50580 $Y=-5
.ENDS
***************************************
.SUBCKT pfet_03v3_I08 1 2 3
** N=3 EP=3 IP=0 FDC=1
XM0 2 3 1 1 pfet_03v3 L=5.6e-07 W=4.2e-07 AD=3.96e-13 AS=3.96e-13 PD=2.68e-06 PS=2.68e-06 NRD=0.488889 NRS=0.488889 m=1 nf=1 $X=0 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nfet_03v3_I15 1 2 3
** N=3 EP=3 IP=0 FDC=1
XM0 2 3 1 1 nfet_03v3 L=5.6e-07 W=2.8e-07 AD=2.64e-13 AS=2.64e-13 PD=2.08e-06 PS=2.08e-06 NRD=0.733333 NRS=0.733333 m=1 nf=1 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pmos_1p2$$48624684
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$47815724
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_28
** N=10 EP=0 IP=12 FDC=0
.ENDS
***************************************
.SUBCKT ICV_29
** N=15 EP=0 IP=20 FDC=0
.ENDS
***************************************
.SUBCKT ICV_30 1 2 3 4 9 11 14 16
** N=16 EP=8 IP=24 FDC=20
*.SEEDPROM
XM0 1 12 10 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=8060 $D=8
XM1 1 15 13 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=9340 $D=8
XM2 12 10 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=8060 $D=8
XM3 15 13 1 1 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=9340 $D=8
X4 3 4 2 2 2 9 11 10 12 018SRAM_cell1_2x $T=0 0 0 0 $X=-340 $Y=-340
X5 3 4 2 2 2 13 15 14 16 018SRAM_cell1_2x $T=0 9000 0 0 $X=-340 $Y=8660
.ENDS
***************************************
.SUBCKT ICV_31 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26
+ 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49
** N=53 EP=40 IP=82 FDC=220
*.SEEDPROM
XM0 7 51 50 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=17060 $D=8
XM1 7 53 52 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=18340 $D=8
XM2 51 50 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=17060 $D=8
XM3 53 52 7 7 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=18340 $D=8
X4 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 30 31
+ 32 33 34 35 36 37 38 39 40 41 42 43 44 45
+ ICV_14 $T=-3000 0 1 180 $X=-15340 $Y=-340
X7 7 8 25 26 46 47 50 51 ICV_30 $T=0 0 0 0 $X=-340 $Y=-340
X8 7 8 25 26 52 53 48 49 ICV_30 $T=0 18000 0 0 $X=-340 $Y=17660
.ENDS
***************************************
.SUBCKT 018SRAM_cell1_dummy_R
** N=8 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_1
** N=11 EP=0 IP=14 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_2 3 4 8 9 10 11
** N=16 EP=6 IP=22 FDC=4
*.SEEDPROM
XM0 4 4 8 4 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=3560 $D=8
XM1 4 4 10 4 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=4840 $D=8
XM2 9 3 4 4 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=3560 $D=8
XM3 11 3 4 4 pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=4840 $D=8
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 10 12 14 15
** N=19 EP=8 IP=26 FDC=16
*.SEEDPROM
XM0 1 3 16 3 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=3180 $Y=7970 $D=2
XM1 18 3 1 3 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=3180 $Y=9260 $D=2
XM2 3 4 16 3 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=3630 $Y=6340 $D=2
XM3 3 4 18 3 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=3630 $Y=10710 $D=2
XM4 17 3 3 3 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=4770 $Y=6340 $D=2
XM5 19 3 3 3 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=4770 $Y=10710 $D=2
XM6 2 3 17 3 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=5220 $Y=7970 $D=2
XM7 19 3 2 3 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=5220 $Y=9260 $D=2
X8 3 4 10 12 16 17 ICV_2 $T=0 0 0 0 $X=-340 $Y=-340
X9 3 4 18 19 14 15 ICV_2 $T=0 9000 0 0 $X=-340 $Y=8660
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 14 16 18 19
** N=23 EP=8 IP=30 FDC=40
*.SEEDPROM
XM0 1 3 20 3 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=3180 $Y=16970 $D=2
XM1 22 3 1 3 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=3180 $Y=18260 $D=2
XM2 3 4 20 3 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=3630 $Y=15340 $D=2
XM3 3 4 22 3 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=3630 $Y=19710 $D=2
XM4 21 3 3 3 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=4770 $Y=15340 $D=2
XM5 23 3 3 3 nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=4770 $Y=19710 $D=2
XM6 2 3 21 3 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=5220 $Y=16970 $D=2
XM7 23 3 2 3 nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=5220 $Y=18260 $D=2
X8 1 2 3 4 14 16 20 21 ICV_3 $T=0 0 0 0 $X=-340 $Y=-340
X9 1 2 3 4 22 23 18 19 ICV_3 $T=0 18000 0 0 $X=-340 $Y=17660
.ENDS
***************************************
.SUBCKT gf180mcu_ocd_ip_sram__sram512x8m8wm1 A[8] A[7] A[6] A[5] A[4] A[3] A[2]
+ A[1] A[0] CEN CLK D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] GWEN Q[7] Q[6]
+ Q[5] Q[4] Q[3] Q[2] Q[1] Q[0] VDD VSS WEN[7] WEN[6] WEN[5] WEN[4] WEN[3]
+ WEN[2] WEN[1] WEN[0]
** N=24897 EP=38 IP=4916 FDC=29933
XM0 23498 VSS 703 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=120390 $Y=176390 $D=2
XM1 703 VSS 23500 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=120390 $Y=472100 $D=2
XM2 VSS 23497 23498 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=120840 $Y=177840 $D=2
XM3 VSS 23499 23500 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=120840 $Y=470470 $D=2
XM4 23497 23498 VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=121980 $Y=177840 $D=2
XM5 23499 23500 VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=121980 $Y=470470 $D=2
XM6 23497 VSS 702 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=122430 $Y=176390 $D=2
XM7 702 VSS 23499 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=122430 $Y=472100 $D=2
XM8 VSS 24106 23202 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=168355 $Y=180895 $D=2
XM9 24106 24042 VSS VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=183295 $D=2
XM10 VSS 24044 24108 VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=213375 $D=2
XM11 VSS 24108 23209 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=214655 $D=2
XM12 VSS 24110 23210 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=216895 $D=2
XM13 24110 24046 VSS VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=219295 $D=2
XM14 VSS 24048 24112 VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=249375 $D=2
XM15 VSS 24112 23217 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=250655 $D=2
XM16 VSS 24114 23218 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=252895 $D=2
XM17 24114 24050 VSS VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=255295 $D=2
XM18 VSS 24052 24116 VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=285375 $D=2
XM19 VSS 24116 23225 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=286655 $D=2
XM20 VSS 24118 23226 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=288895 $D=2
XM21 24118 24054 VSS VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=291295 $D=2
XM22 VSS 24056 24120 VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=321375 $D=2
XM23 VSS 24120 23233 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=322655 $D=2
XM24 VSS 24122 23234 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=324895 $D=2
XM25 24122 24058 VSS VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=327295 $D=2
XM26 VSS 24060 24124 VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=357375 $D=2
XM27 VSS 24124 23241 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=358655 $D=2
XM28 VSS 24126 23242 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=360895 $D=2
XM29 24126 24062 VSS VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=363295 $D=2
XM30 VSS 24064 24128 VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=393375 $D=2
XM31 VSS 24128 23249 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=394655 $D=2
XM32 VSS 24130 23250 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=396895 $D=2
XM33 24130 24066 VSS VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=399295 $D=2
XM34 VSS 24068 24132 VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=429375 $D=2
XM35 VSS 24132 23257 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=430655 $D=2
XM36 VSS 24134 23258 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=168355 $Y=432895 $D=2
XM37 24134 24070 VSS VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=168355 $Y=435295 $D=2
XM38 VSS 24072 24136 VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=168355 $Y=465375 $D=2
XM39 VSS 24136 23265 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=168355 $Y=466655 $D=2
XM40 24042 24043 VSS VSS nfet_03v3 L=2.8e-07 W=1.025e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=198635 $Y=180895 $D=2
XM41 VSS 24045 24044 VSS nfet_03v3 L=2.8e-07 W=1.025e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=198635 $Y=215775 $D=2
XM42 24046 24047 VSS VSS nfet_03v3 L=2.8e-07 W=1.025e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=198635 $Y=216895 $D=2
XM43 VSS 24049 24048 VSS nfet_03v3 L=2.8e-07 W=1.025e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=198635 $Y=251775 $D=2
XM44 24050 24051 VSS VSS nfet_03v3 L=2.8e-07 W=1.025e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=198635 $Y=252895 $D=2
XM45 VSS 24053 24052 VSS nfet_03v3 L=2.8e-07 W=1.025e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=198635 $Y=287775 $D=2
XM46 24054 24055 VSS VSS nfet_03v3 L=2.8e-07 W=1.025e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=198635 $Y=288895 $D=2
XM47 VSS 24057 24056 VSS nfet_03v3 L=2.8e-07 W=1.025e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=198635 $Y=323775 $D=2
XM48 24058 24059 VSS VSS nfet_03v3 L=2.8e-07 W=1.025e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=198635 $Y=324895 $D=2
XM49 VSS 24061 24060 VSS nfet_03v3 L=2.8e-07 W=1.025e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=198635 $Y=359775 $D=2
XM50 24062 24063 VSS VSS nfet_03v3 L=2.8e-07 W=1.025e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=198635 $Y=360895 $D=2
XM51 VSS 24065 24064 VSS nfet_03v3 L=2.8e-07 W=1.025e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=198635 $Y=395775 $D=2
XM52 24066 24067 VSS VSS nfet_03v3 L=2.8e-07 W=1.025e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=198635 $Y=396895 $D=2
XM53 VSS 24069 24068 VSS nfet_03v3 L=2.8e-07 W=1.025e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=198635 $Y=431775 $D=2
XM54 24070 24071 VSS VSS nfet_03v3 L=2.8e-07 W=1.025e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=198635 $Y=432895 $D=2
XM55 VSS 24073 24072 VSS nfet_03v3 L=2.8e-07 W=1.025e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=198635 $Y=467775 $D=2
XM56 2 VDD 1 VSS nfet_03v3 L=2.8e-07 W=3.075e-06 AD=2.8996e-12 AS=2.8996e-12 PD=1.406e-05 PS=1.406e-05 NRD=0.0667678 NRS=0.0667678 m=1 nf=1 $X=204815 $Y=471000 $D=2
XM57 24707 1040 VSS VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=7.32375e-13 AS=2.079e-12 PD=3.615e-06 PS=7.62e-06 NRD=0.0738095 NRS=0.209524 m=1 nf=1 $X=218475 $Y=180950 $D=2
XM58 24706 1044 24707 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=182015 $D=2
XM59 24043 1052 24706 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=183135 $D=2
XM60 24708 1045 24045 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=213535 $D=2
XM61 24709 1044 24708 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=214655 $D=2
XM62 VSS 1040 24709 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=218475 $Y=215720 $D=2
XM63 24711 1040 VSS VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=218475 $Y=216950 $D=2
XM64 24710 1043 24711 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=218015 $D=2
XM65 24047 1052 24710 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=219135 $D=2
XM66 24712 1045 24049 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=249535 $D=2
XM67 24713 1043 24712 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=250655 $D=2
XM68 VSS 1040 24713 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=218475 $Y=251720 $D=2
XM69 24715 1040 VSS VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=218475 $Y=252950 $D=2
XM70 24714 1042 24715 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=254015 $D=2
XM71 24051 1052 24714 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=255135 $D=2
XM72 24716 1045 24053 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=285535 $D=2
XM73 24717 1042 24716 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=286655 $D=2
XM74 VSS 1040 24717 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=218475 $Y=287720 $D=2
XM75 24719 1040 VSS VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=218475 $Y=288950 $D=2
XM76 24718 1041 24719 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=290015 $D=2
XM77 24055 1052 24718 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=291135 $D=2
XM78 24720 1045 24057 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=321535 $D=2
XM79 24721 1041 24720 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=322655 $D=2
XM80 VSS 1040 24721 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=218475 $Y=323720 $D=2
XM81 24723 1038 VSS VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=218475 $Y=324950 $D=2
XM82 24722 1044 24723 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=326015 $D=2
XM83 24059 1052 24722 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=327135 $D=2
XM84 24724 1045 24061 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=357535 $D=2
XM85 24725 1044 24724 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=358655 $D=2
XM86 VSS 1038 24725 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=218475 $Y=359720 $D=2
XM87 24727 1038 VSS VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=218475 $Y=360950 $D=2
XM88 24726 1043 24727 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=362015 $D=2
XM89 24063 1052 24726 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=363135 $D=2
XM90 24728 1045 24065 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=393535 $D=2
XM91 24729 1043 24728 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=394655 $D=2
XM92 VSS 1038 24729 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=218475 $Y=395720 $D=2
XM93 24731 1038 VSS VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=218475 $Y=396950 $D=2
XM94 24730 1042 24731 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=398015 $D=2
XM95 24067 1052 24730 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=399135 $D=2
XM96 24732 1045 24069 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=429535 $D=2
XM97 24733 1042 24732 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=430655 $D=2
XM98 VSS 1038 24733 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=218475 $Y=431720 $D=2
XM99 24735 1038 VSS VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=218475 $Y=432950 $D=2
XM100 24734 1041 24735 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=218475 $Y=434015 $D=2
XM101 24071 1052 24734 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=218475 $Y=435135 $D=2
XM102 24736 1045 24073 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=218475 $Y=465535 $D=2
XM103 24737 1041 24736 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=218475 $Y=466655 $D=2
XM104 VSS 1038 24737 VSS nfet_03v3 L=2.8e-07 W=1.47e-06 AD=2.079e-12 AS=7.32375e-13 PD=7.62e-06 PS=3.615e-06 NRD=0.209524 NRS=0.0738095 m=1 nf=1 $X=218475 $Y=467720 $D=2
XM105 VSS 1 1000 VSS nfet_03v3 L=2.8e-07 W=6.3e-07 AD=3.536e-13 AS=5.984e-13 PD=1.88e-06 PS=3.6e-06 NRD=0.191176 NRS=0.323529 m=1 nf=1 $X=233770 $Y=54135 $D=2
XM106 1000 CLK VSS VSS nfet_03v3 L=2.8e-07 W=6.3e-07 AD=5.984e-13 AS=3.536e-13 PD=3.6e-06 PS=1.88e-06 NRD=0.323529 NRS=0.191176 m=1 nf=1 $X=234890 $Y=54135 $D=2
XM107 616 619 VSS VSS nfet_03v3 L=2.8e-07 W=2.115e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=242235 $Y=54135 $D=2
XM108 281 1006 VSS VSS nfet_03v3 L=4.65e-07 W=2.8e-07 AD=2.64e-13 AS=2.64e-13 PD=2.08e-06 PS=2.08e-06 NRD=0.733333 NRS=0.733333 m=1 nf=1 $X=243265 $Y=46010 $D=2
XM109 CEN 1000 619 VSS nfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=245925 $Y=54135 $D=2
XM110 250 468 VSS VSS nfet_03v3 L=2.8e-07 W=2.329e-05 AD=1.47704e-11 AS=1.47704e-11 PD=6.284e-05 PS=6.284e-05 NRD=0.148297 NRS=0.148297 m=1 nf=5 $X=241995 $Y=72320 $D=2
XM111 317 281 VSS VSS nfet_03v3 L=2.8e-07 W=3.5e-07 AD=3.3e-13 AS=3.3e-13 PD=2.38e-06 PS=2.38e-06 NRD=0.586667 NRS=0.586667 m=1 nf=1 $X=246495 $Y=46075 $D=2
XM112 354 317 VSS VSS nfet_03v3 L=2.8e-07 W=1.405e-06 AD=1.3288e-12 AS=1.3288e-12 PD=6.92e-06 PS=6.92e-06 NRD=0.145695 NRS=0.145695 m=1 nf=1 $X=249065 $Y=46070 $D=2
XM113 24027 354 VSS VSS nfet_03v3 L=2.8e-07 W=1.058e-05 AD=5.8968e-12 AS=1.34946e-11 PD=2.32e-05 PS=4.655e-05 NRD=0.0114638 NRS=0.0262346 m=1 nf=1 $X=256125 $Y=28435 $D=2
XM114 VSS 24107 23266 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=252270 $Y=180895 $D=2
XM115 24107 24042 VSS VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=183295 $D=2
XM116 VSS 24044 24109 VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=213375 $D=2
XM117 VSS 24109 23273 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=214655 $D=2
XM118 VSS 24111 23274 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=216895 $D=2
XM119 24111 24046 VSS VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=219295 $D=2
XM120 VSS 24048 24113 VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=249375 $D=2
XM121 VSS 24113 23281 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=250655 $D=2
XM122 VSS 24115 23282 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=252895 $D=2
XM123 24115 24050 VSS VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=255295 $D=2
XM124 VSS 24052 24117 VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=285375 $D=2
XM125 VSS 24117 23289 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=286655 $D=2
XM126 VSS 24119 23290 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=288895 $D=2
XM127 24119 24054 VSS VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=291295 $D=2
XM128 VSS 24056 24121 VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=321375 $D=2
XM129 VSS 24121 23297 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=322655 $D=2
XM130 VSS 24123 23298 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=324895 $D=2
XM131 24123 24058 VSS VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=327295 $D=2
XM132 VSS 24060 24125 VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=357375 $D=2
XM133 VSS 24125 23305 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=358655 $D=2
XM134 VSS 24127 23306 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=360895 $D=2
XM135 24127 24062 VSS VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=363295 $D=2
XM136 VSS 24064 24129 VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=393375 $D=2
XM137 VSS 24129 23313 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=394655 $D=2
XM138 VSS 24131 23314 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=396895 $D=2
XM139 24131 24066 VSS VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=399295 $D=2
XM140 VSS 24068 24133 VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=429375 $D=2
XM141 VSS 24133 23321 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=430655 $D=2
XM142 VSS 24135 23322 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=252270 $Y=432895 $D=2
XM143 24135 24070 VSS VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=252270 $Y=435295 $D=2
XM144 VSS 24072 24137 VSS nfet_03v3 L=2.8e-07 W=2.33e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=252270 $Y=465375 $D=2
XM145 VSS 24137 23329 VSS nfet_03v3 L=2.8e-07 W=4.665e-06 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=252270 $Y=466655 $D=2
XM146 24028 CLK 24027 VSS nfet_03v3 L=2.8e-07 W=1.058e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=257245 $Y=28435 $D=2
XM147 445 616 24028 VSS nfet_03v3 L=2.8e-07 W=1.058e-05 AD=1.33812e-11 AS=5.8968e-12 PD=4.654e-05 PS=2.32e-05 NRD=0.0260141 NRS=0.0114638 m=1 nf=1 $X=258365 $Y=28435 $D=2
XM148 24029 495 VSS VSS nfet_03v3 L=2.8e-07 W=8.465e-06 AD=4.7177e-12 AS=1.07963e-11 PD=1.8665e-05 PS=3.748e-05 NRD=0.014329 NRS=0.0327914 m=1 nf=1 $X=262120 $Y=29545 $D=2
XM149 468 445 24029 VSS nfet_03v3 L=2.8e-07 W=8.465e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=263240 $Y=29545 $D=2
XM150 24030 445 468 VSS nfet_03v3 L=2.8e-07 W=8.465e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=264360 $Y=29545 $D=2
XM151 VSS 495 24030 VSS nfet_03v3 L=2.8e-07 W=8.465e-06 AD=1.07055e-11 AS=4.7177e-12 PD=3.747e-05 PS=1.8665e-05 NRD=0.0325158 NRS=0.014329 m=1 nf=1 $X=265480 $Y=29545 $D=2
XM152 24031 468 VSS VSS nfet_03v3 L=2.8e-07 W=2.115e-06 AD=1.16905e-12 AS=2.7013e-12 PD=5.055e-06 PS=1.027e-05 NRD=0.0567181 NRS=0.131057 m=1 nf=1 $X=268545 $Y=43150 $D=2
XM153 495 607 24031 VSS nfet_03v3 L=2.8e-07 W=2.115e-06 AD=2.27e-14 AS=-2.27e-14 PD=1e-08 PS=-1e-08 NRD=0.00110132 NRS=-0.00110132 m=1 nf=1 $X=269660 $Y=43150 $D=2
XM154 24032 607 495 VSS nfet_03v3 L=2.8e-07 W=2.115e-06 AD=-2.27e-14 AS=2.27e-14 PD=-1e-08 PS=1e-08 NRD=-0.00110132 NRS=0.00110132 m=1 nf=1 $X=270785 $Y=43150 $D=2
XM155 VSS 468 24032 VSS nfet_03v3 L=2.8e-07 W=2.115e-06 AD=2.7013e-12 AS=1.16905e-12 PD=1.027e-05 PS=5.055e-06 NRD=0.131057 NRS=0.0567181 m=1 nf=1 $X=271900 $Y=43150 $D=2
XM156 1 250 VSS VSS nfet_03v3 L=2.8e-07 W=6.87e-05 AD=3.8324e-11 AS=4.09772e-11 PD=0.0001578 PS=0.00017326 NRD=0.705563 NRS=0.75441 m=1 nf=20 $X=253180 $Y=76320 $D=2
XM157 23502 VSS 705 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=304270 $Y=176390 $D=2
XM158 705 VSS 23504 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=304270 $Y=472100 $D=2
XM159 VSS 23501 23502 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=304720 $Y=177840 $D=2
XM160 VSS 23503 23504 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=304720 $Y=470470 $D=2
XM161 23501 23502 VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=305860 $Y=177840 $D=2
XM162 23503 23504 VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=305860 $Y=470470 $D=2
XM163 23501 VSS 704 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=306310 $Y=176390 $D=2
XM164 704 VSS 23503 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=306310 $Y=472100 $D=2
XM165 24074 VSS 614 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=418270 $Y=176390 $D=2
XM166 614 VSS 24076 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=211100 $D=2
XM167 24078 VSS 614 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=212390 $D=2
XM168 614 VSS 24080 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=247100 $D=2
XM169 24082 VSS 614 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=248390 $D=2
XM170 614 VSS 24084 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=283100 $D=2
XM171 24086 VSS 614 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=284390 $D=2
XM172 614 VSS 24088 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=319100 $D=2
XM173 24090 VSS 614 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=320390 $D=2
XM174 614 VSS 24092 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=355100 $D=2
XM175 24094 VSS 614 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=356390 $D=2
XM176 614 VSS 24096 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=391100 $D=2
XM177 24098 VSS 614 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=392390 $D=2
XM178 614 VSS 24100 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=427100 $D=2
XM179 24102 VSS 614 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=428390 $D=2
XM180 614 1002 24104 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=463100 $D=2
XM181 23859 1002 614 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=464390 $D=2
XM182 614 1002 23857 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=418270 $Y=472100 $D=2
XM183 VSS VDD 24074 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=177840 $D=2
XM184 VSS VDD 24076 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=209470 $D=2
XM185 VSS VDD 24078 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=213840 $D=2
XM186 VSS VDD 24080 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=245470 $D=2
XM187 VSS VDD 24082 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=249840 $D=2
XM188 VSS VDD 24084 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=281470 $D=2
XM189 VSS VDD 24086 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=285840 $D=2
XM190 VSS VDD 24088 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=317470 $D=2
XM191 VSS VDD 24090 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=321840 $D=2
XM192 VSS VDD 24092 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=353470 $D=2
XM193 VSS VDD 24094 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=357840 $D=2
XM194 VSS VDD 24096 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=389470 $D=2
XM195 VSS VDD 24098 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=393840 $D=2
XM196 VSS VDD 24100 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=425470 $D=2
XM197 VSS VDD 24102 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=429840 $D=2
XM198 VSS VDD 24104 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=461470 $D=2
XM199 VSS VDD 23859 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=465840 $D=2
XM200 VSS VDD 23857 VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=470470 $D=2
XM201 24075 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=177840 $D=2
XM202 24077 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=209470 $D=2
XM203 24079 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=213840 $D=2
XM204 24081 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=245470 $D=2
XM205 24083 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=249840 $D=2
XM206 24085 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=281470 $D=2
XM207 24087 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=285840 $D=2
XM208 24089 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=317470 $D=2
XM209 24091 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=321840 $D=2
XM210 24093 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=353470 $D=2
XM211 24095 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=357840 $D=2
XM212 24097 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=389470 $D=2
XM213 24099 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=393840 $D=2
XM214 24101 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=425470 $D=2
XM215 24103 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=429840 $D=2
XM216 24105 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=461470 $D=2
XM217 23860 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=465840 $D=2
XM218 23858 VSS VSS VSS nfet_03v3 L=2.8e-07 W=4.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=470470 $D=2
XM219 606 614 VSS VSS nfet_03v3 L=2.8e-07 W=1.285e-06 AD=7.176e-13 AS=1.2144e-12 PD=3.8e-06 PS=7.28e-06 NRD=0.376812 NRS=0.637681 m=1 nf=2 $X=418770 $Y=94540 $D=2
XM220 607 606 VSS VSS nfet_03v3 L=2.8e-07 W=7.93e-06 AD=4.42e-12 AS=7.48e-12 PD=1.804e-05 PS=3.576e-05 NRD=0.0611765 NRS=0.103529 m=1 nf=2 $X=418790 $Y=79115 $D=2
XM221 613 VDD VSS VSS nfet_03v3 L=2.8e-07 W=5.3e-07 AD=2.964e-13 AS=5.016e-13 PD=2.18e-06 PS=4.04e-06 NRD=0.912281 NRS=1.54386 m=1 nf=2 $X=419015 $Y=110805 $D=2
XM222 24075 VSS 615 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=420310 $Y=176390 $D=2
XM223 615 VSS 24077 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=211100 $D=2
XM224 24079 VSS 615 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=212390 $D=2
XM225 615 VSS 24081 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=247100 $D=2
XM226 24083 VSS 615 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=248390 $D=2
XM227 615 VSS 24085 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=283100 $D=2
XM228 24087 VSS 615 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=284390 $D=2
XM229 615 VSS 24089 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=319100 $D=2
XM230 24091 VSS 615 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=320390 $D=2
XM231 615 VSS 24093 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=355100 $D=2
XM232 24095 VSS 615 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=356390 $D=2
XM233 615 VSS 24097 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=391100 $D=2
XM234 24099 VSS 615 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=392390 $D=2
XM235 615 VSS 24101 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=427100 $D=2
XM236 24103 VSS 615 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=428390 $D=2
XM237 615 1002 24105 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=463100 $D=2
XM238 23860 1002 615 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=464390 $D=2
XM239 615 1002 23858 VSS nfet_03v3 L=3.6e-07 W=2.8e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=420310 $Y=472100 $D=2
XM240 VDD 23446 23448 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=179690 $D=8
XM241 VDD 24167 24166 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=180970 $D=8
XM242 VDD 24175 24174 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=323690 $D=8
XM243 VDD 24183 24182 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=324970 $D=8
XM244 VDD 24191 24190 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=467690 $D=8
XM245 VDD 23534 23536 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=468970 $D=8
XM246 23446 23448 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=179690 $D=8
XM247 24167 24166 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=180970 $D=8
XM248 24175 24174 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=323690 $D=8
XM249 24183 24182 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=324970 $D=8
XM250 24191 24190 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=467690 $D=8
XM251 23534 23536 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=468970 $D=8
XM252 23915 23198 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=13620 $Y=160970 $D=8
XM253 23916 23198 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=13620 $Y=164845 $D=8
XM254 24138 23885 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=13835 $Y=112830 $D=8
XM255 VDD 23442 23444 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=179690 $D=8
XM256 VDD 24169 24168 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=180970 $D=8
XM257 VDD 24177 24176 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=323690 $D=8
XM258 VDD 24185 24184 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=324970 $D=8
XM259 VDD 24193 24192 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=467690 $D=8
XM260 VDD 23530 23532 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=468970 $D=8
XM261 23442 23444 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=179690 $D=8
XM262 24169 24168 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=180970 $D=8
XM263 24177 24176 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=323690 $D=8
XM264 24185 24184 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=324970 $D=8
XM265 24193 24192 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=467690 $D=8
XM266 23530 23532 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=468970 $D=8
XM267 24139 23884 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=16365 $Y=112830 $D=8
XM268 23918 23198 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=16720 $Y=160970 $D=8
XM269 23917 23198 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=16720 $Y=164845 $D=8
XM270 VDD 23438 23440 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=179690 $D=8
XM271 VDD 24171 24170 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=180970 $D=8
XM272 VDD 24179 24178 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=323690 $D=8
XM273 VDD 24187 24186 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=324970 $D=8
XM274 VDD 24195 24194 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=467690 $D=8
XM275 VDD 23526 23528 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=468970 $D=8
XM276 23438 23440 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=179690 $D=8
XM277 24171 24170 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=180970 $D=8
XM278 24179 24178 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=323690 $D=8
XM279 24187 24186 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=324970 $D=8
XM280 24195 24194 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=467690 $D=8
XM281 23526 23528 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=468970 $D=8
XM282 23919 23198 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=19815 $Y=160970 $D=8
XM283 23920 23198 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=19815 $Y=164845 $D=8
XM284 24140 23883 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=20030 $Y=112830 $D=8
XM285 VDD 23434 23436 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=179690 $D=8
XM286 VDD 24173 24172 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=180970 $D=8
XM287 VDD 24181 24180 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=323690 $D=8
XM288 VDD 24189 24188 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=324970 $D=8
XM289 VDD 24197 24196 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=467690 $D=8
XM290 VDD 23522 23524 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=468970 $D=8
XM291 23434 23436 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=179690 $D=8
XM292 24173 24172 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=180970 $D=8
XM293 24181 24180 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=323690 $D=8
XM294 24189 24188 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=324970 $D=8
XM295 24197 24196 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=467690 $D=8
XM296 23522 23524 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=468970 $D=8
XM297 24141 23882 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=22560 $Y=112830 $D=8
XM298 23922 23198 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=22915 $Y=160970 $D=8
XM299 23921 23198 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=22915 $Y=164845 $D=8
XM300 VDD 23342 23344 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=179690 $D=8
XM301 VDD 24263 24262 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=180970 $D=8
XM302 VDD 24287 24286 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=323690 $D=8
XM303 VDD 24311 24310 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=324970 $D=8
XM304 VDD 24335 24334 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=467690 $D=8
XM305 VDD 23518 23520 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=468970 $D=8
XM306 23342 23344 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=179690 $D=8
XM307 24263 24262 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=180970 $D=8
XM308 24287 24286 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=323690 $D=8
XM309 24311 24310 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=324970 $D=8
XM310 24335 24334 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=467690 $D=8
XM311 23518 23520 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=468970 $D=8
XM312 23923 23198 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=26005 $Y=160970 $D=8
XM313 23924 23198 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=26005 $Y=164845 $D=8
XM314 24142 23881 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=26220 $Y=112830 $D=8
XM315 VDD 23338 23340 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=179690 $D=8
XM316 VDD 24265 24264 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=180970 $D=8
XM317 VDD 24289 24288 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=323690 $D=8
XM318 VDD 24313 24312 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=324970 $D=8
XM319 VDD 24337 24336 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=467690 $D=8
XM320 VDD 23514 23516 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=468970 $D=8
XM321 23338 23340 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=179690 $D=8
XM322 24265 24264 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=180970 $D=8
XM323 24289 24288 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=323690 $D=8
XM324 24313 24312 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=324970 $D=8
XM325 24337 24336 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=467690 $D=8
XM326 23514 23516 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=468970 $D=8
XM327 24143 23880 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=28750 $Y=112830 $D=8
XM328 23926 23198 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=29105 $Y=160970 $D=8
XM329 23925 23198 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=29105 $Y=164845 $D=8
XM330 VDD 23350 23352 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=179690 $D=8
XM331 VDD 24267 24266 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=180970 $D=8
XM332 VDD 24291 24290 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=323690 $D=8
XM333 VDD 24315 24314 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=324970 $D=8
XM334 VDD 24339 24338 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=467690 $D=8
XM335 VDD 23510 23512 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=468970 $D=8
XM336 23350 23352 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=179690 $D=8
XM337 24267 24266 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=180970 $D=8
XM338 24291 24290 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=323690 $D=8
XM339 24315 24314 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=324970 $D=8
XM340 24339 24338 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=467690 $D=8
XM341 23510 23512 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=468970 $D=8
XM342 23927 23198 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=32200 $Y=160970 $D=8
XM343 23928 23198 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=32200 $Y=164845 $D=8
XM344 24144 23879 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=32415 $Y=112830 $D=8
XM345 VDD 23346 23348 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=179690 $D=8
XM346 VDD 24269 24268 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=180970 $D=8
XM347 VDD 24293 24292 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=323690 $D=8
XM348 VDD 24317 24316 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=324970 $D=8
XM349 VDD 24341 24340 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=467690 $D=8
XM350 VDD 23506 23508 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=468970 $D=8
XM351 23346 23348 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=179690 $D=8
XM352 24269 24268 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=180970 $D=8
XM353 24293 24292 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=323690 $D=8
XM354 24317 24316 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=324970 $D=8
XM355 24341 24340 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=467690 $D=8
XM356 23506 23508 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=468970 $D=8
XM357 24034 23878 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=34945 $Y=112830 $D=8
XM358 1064 23198 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=35120 $Y=160970 $D=8
XM359 1065 23198 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=35120 $Y=164845 $D=8
XM360 1076 1074 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=38575 $Y=160970 $D=8
XM361 1077 1074 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=38575 $Y=164845 $D=8
XM362 VDD 23566 23568 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=179690 $D=8
XM363 VDD 24284 24285 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=180970 $D=8
XM364 VDD 24308 24309 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=323690 $D=8
XM365 VDD 24332 24333 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=324970 $D=8
XM366 VDD 24356 24357 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=467690 $D=8
XM367 VDD 23598 23600 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=468970 $D=8
XM368 24038 23885 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=38620 $Y=112830 $D=8
XM369 23566 23568 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=179690 $D=8
XM370 24284 24285 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=180970 $D=8
XM371 24308 24309 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=323690 $D=8
XM372 24332 24333 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=324970 $D=8
XM373 24356 24357 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=467690 $D=8
XM374 23598 23600 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=468970 $D=8
XM375 24652 23884 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=41145 $Y=112830 $D=8
XM376 23983 1074 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=41500 $Y=160970 $D=8
XM377 23984 1074 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=41500 $Y=164845 $D=8
XM378 VDD 23562 23564 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=179690 $D=8
XM379 VDD 24282 24283 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=180970 $D=8
XM380 VDD 24306 24307 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=323690 $D=8
XM381 VDD 24330 24331 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=324970 $D=8
XM382 VDD 24354 24355 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=467690 $D=8
XM383 VDD 23594 23596 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=468970 $D=8
XM384 23562 23564 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=179690 $D=8
XM385 24282 24283 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=180970 $D=8
XM386 24306 24307 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=323690 $D=8
XM387 24330 24331 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=324970 $D=8
XM388 24354 24355 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=467690 $D=8
XM389 23594 23596 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=468970 $D=8
XM390 23982 1074 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=44595 $Y=160970 $D=8
XM391 23981 1074 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=44595 $Y=164845 $D=8
XM392 VDD 23558 23560 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=179690 $D=8
XM393 VDD 24280 24281 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=180970 $D=8
XM394 VDD 24304 24305 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=323690 $D=8
XM395 VDD 24328 24329 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=324970 $D=8
XM396 VDD 24352 24353 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=467690 $D=8
XM397 VDD 23590 23592 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=468970 $D=8
XM398 24651 23883 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=44810 $Y=112830 $D=8
XM399 23558 23560 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=179690 $D=8
XM400 24280 24281 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=180970 $D=8
XM401 24304 24305 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=323690 $D=8
XM402 24328 24329 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=324970 $D=8
XM403 24352 24353 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=467690 $D=8
XM404 23590 23592 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=468970 $D=8
XM405 24650 23882 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=47340 $Y=112830 $D=8
XM406 23979 1074 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=47695 $Y=160970 $D=8
XM407 23980 1074 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=47695 $Y=164845 $D=8
XM408 VDD 23554 23556 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=179690 $D=8
XM409 VDD 24278 24279 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=180970 $D=8
XM410 VDD 24302 24303 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=323690 $D=8
XM411 VDD 24326 24327 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=324970 $D=8
XM412 VDD 24350 24351 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=467690 $D=8
XM413 VDD 23586 23588 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=468970 $D=8
XM414 23554 23556 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=179690 $D=8
XM415 24278 24279 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=180970 $D=8
XM416 24302 24303 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=323690 $D=8
XM417 24326 24327 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=324970 $D=8
XM418 24350 24351 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=467690 $D=8
XM419 23586 23588 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=468970 $D=8
XM420 VDD 23550 23552 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=179690 $D=8
XM421 VDD 24276 24277 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=180970 $D=8
XM422 VDD 24300 24301 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=323690 $D=8
XM423 VDD 24324 24325 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=324970 $D=8
XM424 VDD 24348 24349 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=467690 $D=8
XM425 VDD 23582 23584 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=468970 $D=8
XM426 23978 1074 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=50785 $Y=160970 $D=8
XM427 23977 1074 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=50785 $Y=164845 $D=8
XM428 24649 23881 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=51000 $Y=112830 $D=8
XM429 23550 23552 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=179690 $D=8
XM430 24276 24277 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=180970 $D=8
XM431 24300 24301 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=323690 $D=8
XM432 24324 24325 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=324970 $D=8
XM433 24348 24349 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=467690 $D=8
XM434 23582 23584 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=468970 $D=8
XM435 24648 23880 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=53530 $Y=112830 $D=8
XM436 VDD 23546 23548 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=179690 $D=8
XM437 VDD 24274 24275 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=180970 $D=8
XM438 VDD 24298 24299 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=323690 $D=8
XM439 VDD 24322 24323 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=324970 $D=8
XM440 VDD 24346 24347 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=467690 $D=8
XM441 VDD 23578 23580 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=468970 $D=8
XM442 23975 1074 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=53885 $Y=160970 $D=8
XM443 23976 1074 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=53885 $Y=164845 $D=8
XM444 23546 23548 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=179690 $D=8
XM445 24274 24275 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=180970 $D=8
XM446 24298 24299 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=323690 $D=8
XM447 24322 24323 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=324970 $D=8
XM448 24346 24347 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=467690 $D=8
XM449 23578 23580 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=468970 $D=8
XM450 VDD 23542 23544 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=179690 $D=8
XM451 VDD 24272 24273 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=180970 $D=8
XM452 VDD 24296 24297 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=323690 $D=8
XM453 VDD 24320 24321 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=324970 $D=8
XM454 VDD 24344 24345 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=467690 $D=8
XM455 VDD 23574 23576 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=468970 $D=8
XM456 23974 1074 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=56980 $Y=160970 $D=8
XM457 23973 1074 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=56980 $Y=164845 $D=8
XM458 24647 23879 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=57195 $Y=112830 $D=8
XM459 23542 23544 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=179690 $D=8
XM460 24272 24273 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=180970 $D=8
XM461 24296 24297 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=323690 $D=8
XM462 24320 24321 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=324970 $D=8
XM463 24344 24345 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=467690 $D=8
XM464 23574 23576 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=468970 $D=8
XM465 VDD 23538 23540 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=179690 $D=8
XM466 VDD 24270 24271 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=180970 $D=8
XM467 VDD 24294 24295 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=323690 $D=8
XM468 VDD 24318 24319 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=324970 $D=8
XM469 VDD 24342 24343 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=467690 $D=8
XM470 VDD 23570 23572 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=468970 $D=8
XM471 24646 23878 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=59725 $Y=112830 $D=8
XM472 23971 1074 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=60080 $Y=160970 $D=8
XM473 23972 1074 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=60080 $Y=164845 $D=8
XM474 23538 23540 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=179690 $D=8
XM475 24270 24271 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=180970 $D=8
XM476 24294 24295 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=323690 $D=8
XM477 24318 24319 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=324970 $D=8
XM478 24342 24343 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=467690 $D=8
XM479 23570 23572 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=468970 $D=8
XM480 VDD 23462 23464 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=179690 $D=8
XM481 VDD 24199 24198 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=180970 $D=8
XM482 VDD 24207 24206 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=323690 $D=8
XM483 VDD 24215 24214 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=324970 $D=8
XM484 VDD 24223 24222 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=467690 $D=8
XM485 VDD 23630 23632 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=468970 $D=8
XM486 23462 23464 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=179690 $D=8
XM487 24199 24198 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=180970 $D=8
XM488 24207 24206 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=323690 $D=8
XM489 24215 24214 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=324970 $D=8
XM490 24223 24222 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=467690 $D=8
XM491 23630 23632 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=468970 $D=8
XM492 23929 23199 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=67620 $Y=160970 $D=8
XM493 23930 23199 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=67620 $Y=164845 $D=8
XM494 24145 23885 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=67835 $Y=112830 $D=8
XM495 VDD 23458 23460 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=179690 $D=8
XM496 VDD 24201 24200 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=180970 $D=8
XM497 VDD 24209 24208 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=323690 $D=8
XM498 VDD 24217 24216 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=324970 $D=8
XM499 VDD 24225 24224 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=467690 $D=8
XM500 VDD 23626 23628 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=468970 $D=8
XM501 23458 23460 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=179690 $D=8
XM502 24201 24200 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=180970 $D=8
XM503 24209 24208 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=323690 $D=8
XM504 24217 24216 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=324970 $D=8
XM505 24225 24224 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=467690 $D=8
XM506 23626 23628 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=468970 $D=8
XM507 24146 23884 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=70365 $Y=112830 $D=8
XM508 23932 23199 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=70720 $Y=160970 $D=8
XM509 23931 23199 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=70720 $Y=164845 $D=8
XM510 VDD 23454 23456 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=179690 $D=8
XM511 VDD 24203 24202 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=180970 $D=8
XM512 VDD 24211 24210 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=323690 $D=8
XM513 VDD 24219 24218 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=324970 $D=8
XM514 VDD 24227 24226 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=467690 $D=8
XM515 VDD 23622 23624 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=468970 $D=8
XM516 23454 23456 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=179690 $D=8
XM517 24203 24202 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=180970 $D=8
XM518 24211 24210 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=323690 $D=8
XM519 24219 24218 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=324970 $D=8
XM520 24227 24226 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=467690 $D=8
XM521 23622 23624 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=468970 $D=8
XM522 23933 23199 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=73815 $Y=160970 $D=8
XM523 23934 23199 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=73815 $Y=164845 $D=8
XM524 24147 23883 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=74030 $Y=112830 $D=8
XM525 VDD 23450 23452 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=179690 $D=8
XM526 VDD 24205 24204 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=180970 $D=8
XM527 VDD 24213 24212 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=323690 $D=8
XM528 VDD 24221 24220 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=324970 $D=8
XM529 VDD 24229 24228 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=467690 $D=8
XM530 VDD 23618 23620 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=468970 $D=8
XM531 23450 23452 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=179690 $D=8
XM532 24205 24204 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=180970 $D=8
XM533 24213 24212 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=323690 $D=8
XM534 24221 24220 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=324970 $D=8
XM535 24229 24228 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=467690 $D=8
XM536 23618 23620 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=468970 $D=8
XM537 24148 23882 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=76560 $Y=112830 $D=8
XM538 23936 23199 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=76915 $Y=160970 $D=8
XM539 23935 23199 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=76915 $Y=164845 $D=8
XM540 VDD 23358 23360 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=179690 $D=8
XM541 VDD 24359 24358 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=180970 $D=8
XM542 VDD 24383 24382 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=323690 $D=8
XM543 VDD 24407 24406 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=324970 $D=8
XM544 VDD 24431 24430 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=467690 $D=8
XM545 VDD 23614 23616 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=468970 $D=8
XM546 23358 23360 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=179690 $D=8
XM547 24359 24358 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=180970 $D=8
XM548 24383 24382 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=323690 $D=8
XM549 24407 24406 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=324970 $D=8
XM550 24431 24430 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=467690 $D=8
XM551 23614 23616 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=468970 $D=8
XM552 23937 23199 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=80005 $Y=160970 $D=8
XM553 23938 23199 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=80005 $Y=164845 $D=8
XM554 24149 23881 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=80220 $Y=112830 $D=8
XM555 VDD 23354 23356 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=179690 $D=8
XM556 VDD 24361 24360 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=180970 $D=8
XM557 VDD 24385 24384 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=323690 $D=8
XM558 VDD 24409 24408 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=324970 $D=8
XM559 VDD 24433 24432 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=467690 $D=8
XM560 VDD 23610 23612 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=468970 $D=8
XM561 23354 23356 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=179690 $D=8
XM562 24361 24360 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=180970 $D=8
XM563 24385 24384 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=323690 $D=8
XM564 24409 24408 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=324970 $D=8
XM565 24433 24432 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=467690 $D=8
XM566 23610 23612 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=468970 $D=8
XM567 24150 23880 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=82750 $Y=112830 $D=8
XM568 23940 23199 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=83105 $Y=160970 $D=8
XM569 23939 23199 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=83105 $Y=164845 $D=8
XM570 VDD 23366 23368 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=179690 $D=8
XM571 VDD 24363 24362 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=180970 $D=8
XM572 VDD 24387 24386 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=323690 $D=8
XM573 VDD 24411 24410 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=324970 $D=8
XM574 VDD 24435 24434 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=467690 $D=8
XM575 VDD 23606 23608 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=468970 $D=8
XM576 23366 23368 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=179690 $D=8
XM577 24363 24362 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=180970 $D=8
XM578 24387 24386 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=323690 $D=8
XM579 24411 24410 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=324970 $D=8
XM580 24435 24434 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=467690 $D=8
XM581 23606 23608 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=468970 $D=8
XM582 23941 23199 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=86200 $Y=160970 $D=8
XM583 23942 23199 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=86200 $Y=164845 $D=8
XM584 24151 23879 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=86415 $Y=112830 $D=8
XM585 VDD 23362 23364 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=179690 $D=8
XM586 VDD 24365 24364 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=180970 $D=8
XM587 VDD 24389 24388 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=323690 $D=8
XM588 VDD 24413 24412 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=324970 $D=8
XM589 VDD 24437 24436 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=467690 $D=8
XM590 VDD 23602 23604 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=468970 $D=8
XM591 23362 23364 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=179690 $D=8
XM592 24365 24364 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=180970 $D=8
XM593 24389 24388 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=323690 $D=8
XM594 24413 24412 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=324970 $D=8
XM595 24437 24436 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=467690 $D=8
XM596 23602 23604 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=468970 $D=8
XM597 24035 23878 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=88945 $Y=112830 $D=8
XM598 1066 23199 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=89120 $Y=160970 $D=8
XM599 1067 23199 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=89120 $Y=164845 $D=8
XM600 1079 1078 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=92575 $Y=160970 $D=8
XM601 1080 1078 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=92575 $Y=164845 $D=8
XM602 VDD 23662 23664 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=179690 $D=8
XM603 VDD 24380 24381 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=180970 $D=8
XM604 VDD 24404 24405 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=323690 $D=8
XM605 VDD 24428 24429 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=324970 $D=8
XM606 VDD 24452 24453 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=467690 $D=8
XM607 VDD 23694 23696 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=468970 $D=8
XM608 24039 23885 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=92620 $Y=112830 $D=8
XM609 23662 23664 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=179690 $D=8
XM610 24380 24381 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=180970 $D=8
XM611 24404 24405 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=323690 $D=8
XM612 24428 24429 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=324970 $D=8
XM613 24452 24453 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=467690 $D=8
XM614 23694 23696 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=468970 $D=8
XM615 24659 23884 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=95145 $Y=112830 $D=8
XM616 23997 1078 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=95500 $Y=160970 $D=8
XM617 23998 1078 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=95500 $Y=164845 $D=8
XM618 VDD 23658 23660 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=179690 $D=8
XM619 VDD 24378 24379 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=180970 $D=8
XM620 VDD 24402 24403 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=323690 $D=8
XM621 VDD 24426 24427 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=324970 $D=8
XM622 VDD 24450 24451 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=467690 $D=8
XM623 VDD 23690 23692 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=468970 $D=8
XM624 23658 23660 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=179690 $D=8
XM625 24378 24379 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=180970 $D=8
XM626 24402 24403 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=323690 $D=8
XM627 24426 24427 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=324970 $D=8
XM628 24450 24451 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=467690 $D=8
XM629 23690 23692 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=468970 $D=8
XM630 23996 1078 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=98595 $Y=160970 $D=8
XM631 23995 1078 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=98595 $Y=164845 $D=8
XM632 VDD 23654 23656 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=179690 $D=8
XM633 VDD 24376 24377 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=180970 $D=8
XM634 VDD 24400 24401 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=323690 $D=8
XM635 VDD 24424 24425 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=324970 $D=8
XM636 VDD 24448 24449 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=467690 $D=8
XM637 VDD 23686 23688 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=468970 $D=8
XM638 24658 23883 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=98810 $Y=112830 $D=8
XM639 23654 23656 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=179690 $D=8
XM640 24376 24377 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=180970 $D=8
XM641 24400 24401 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=323690 $D=8
XM642 24424 24425 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=324970 $D=8
XM643 24448 24449 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=467690 $D=8
XM644 23686 23688 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=468970 $D=8
XM645 24657 23882 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=101340 $Y=112830 $D=8
XM646 23993 1078 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=101695 $Y=160970 $D=8
XM647 23994 1078 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=101695 $Y=164845 $D=8
XM648 VDD 23650 23652 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=179690 $D=8
XM649 VDD 24374 24375 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=180970 $D=8
XM650 VDD 24398 24399 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=323690 $D=8
XM651 VDD 24422 24423 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=324970 $D=8
XM652 VDD 24446 24447 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=467690 $D=8
XM653 VDD 23682 23684 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=468970 $D=8
XM654 23650 23652 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=179690 $D=8
XM655 24374 24375 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=180970 $D=8
XM656 24398 24399 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=323690 $D=8
XM657 24422 24423 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=324970 $D=8
XM658 24446 24447 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=467690 $D=8
XM659 23682 23684 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=468970 $D=8
XM660 VDD 23646 23648 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=179690 $D=8
XM661 VDD 24372 24373 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=180970 $D=8
XM662 VDD 24396 24397 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=323690 $D=8
XM663 VDD 24420 24421 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=324970 $D=8
XM664 VDD 24444 24445 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=467690 $D=8
XM665 VDD 23678 23680 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=468970 $D=8
XM666 23992 1078 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=104785 $Y=160970 $D=8
XM667 23991 1078 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=104785 $Y=164845 $D=8
XM668 24656 23881 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=105000 $Y=112830 $D=8
XM669 23646 23648 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=179690 $D=8
XM670 24372 24373 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=180970 $D=8
XM671 24396 24397 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=323690 $D=8
XM672 24420 24421 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=324970 $D=8
XM673 24444 24445 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=467690 $D=8
XM674 23678 23680 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=468970 $D=8
XM675 24655 23880 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=107530 $Y=112830 $D=8
XM676 VDD 23642 23644 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=179690 $D=8
XM677 VDD 24370 24371 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=180970 $D=8
XM678 VDD 24394 24395 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=323690 $D=8
XM679 VDD 24418 24419 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=324970 $D=8
XM680 VDD 24442 24443 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=467690 $D=8
XM681 VDD 23674 23676 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=468970 $D=8
XM682 23989 1078 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=107885 $Y=160970 $D=8
XM683 23990 1078 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=107885 $Y=164845 $D=8
XM684 23642 23644 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=179690 $D=8
XM685 24370 24371 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=180970 $D=8
XM686 24394 24395 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=323690 $D=8
XM687 24418 24419 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=324970 $D=8
XM688 24442 24443 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=467690 $D=8
XM689 23674 23676 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=468970 $D=8
XM690 VDD 23638 23640 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=179690 $D=8
XM691 VDD 24368 24369 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=180970 $D=8
XM692 VDD 24392 24393 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=323690 $D=8
XM693 VDD 24416 24417 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=324970 $D=8
XM694 VDD 24440 24441 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=467690 $D=8
XM695 VDD 23670 23672 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=468970 $D=8
XM696 23988 1078 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=110980 $Y=160970 $D=8
XM697 23987 1078 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=110980 $Y=164845 $D=8
XM698 24654 23879 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=111195 $Y=112830 $D=8
XM699 23638 23640 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=179690 $D=8
XM700 24368 24369 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=180970 $D=8
XM701 24392 24393 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=323690 $D=8
XM702 24416 24417 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=324970 $D=8
XM703 24440 24441 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=467690 $D=8
XM704 23670 23672 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=468970 $D=8
XM705 VDD 23634 23636 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=179690 $D=8
XM706 VDD 24366 24367 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=180970 $D=8
XM707 VDD 24390 24391 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=323690 $D=8
XM708 VDD 24414 24415 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=324970 $D=8
XM709 VDD 24438 24439 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=467690 $D=8
XM710 VDD 23666 23668 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=468970 $D=8
XM711 24653 23878 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=113725 $Y=112830 $D=8
XM712 23985 1078 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=114080 $Y=160970 $D=8
XM713 23986 1078 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=114080 $Y=164845 $D=8
XM714 23634 23636 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=179690 $D=8
XM715 24366 24367 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=180970 $D=8
XM716 24390 24391 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=323690 $D=8
XM717 24414 24415 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=324970 $D=8
XM718 24438 24439 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=467690 $D=8
XM719 23666 23668 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=468970 $D=8
XM720 VDD 23497 23498 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=179690 $D=8
XM721 VDD 24674 24675 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=180970 $D=8
XM722 VDD 24676 24677 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=215690 $D=8
XM723 VDD 24678 24679 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=216970 $D=8
XM724 VDD 24680 24681 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=251690 $D=8
XM725 VDD 24682 24683 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=252970 $D=8
XM726 VDD 24684 24685 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=287690 $D=8
XM727 VDD 24686 24687 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=288970 $D=8
XM728 VDD 24688 24689 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=323690 $D=8
XM729 VDD 24690 24691 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=324970 $D=8
XM730 VDD 24692 24693 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=359690 $D=8
XM731 VDD 24694 24695 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=360970 $D=8
XM732 VDD 24696 24697 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=395690 $D=8
XM733 VDD 24698 24699 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=396970 $D=8
XM734 VDD 24700 24701 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=431690 $D=8
XM735 VDD 24702 24703 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=432970 $D=8
XM736 VDD 24704 24705 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=467690 $D=8
XM737 VDD 23499 23500 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=468970 $D=8
XM738 VDD VSS VDD VDD pfet_03v3 L=1.74e-06 W=3.816e-05 AD=0 AS=6.1309e-11 PD=0 PS=0.000217698 NRD=0 NRS=11.8457 m=1 nf=36 $X=10835 $Y=171065 $D=8
XM739 23497 23498 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=179690 $D=8
XM740 24674 24675 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=180970 $D=8
XM741 24676 24677 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=215690 $D=8
XM742 24678 24679 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=216970 $D=8
XM743 24680 24681 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=251690 $D=8
XM744 24682 24683 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=252970 $D=8
XM745 24684 24685 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=287690 $D=8
XM746 24686 24687 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=288970 $D=8
XM747 24688 24689 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=323690 $D=8
XM748 24690 24691 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=324970 $D=8
XM749 24692 24693 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=359690 $D=8
XM750 24694 24695 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=360970 $D=8
XM751 24696 24697 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=395690 $D=8
XM752 24698 24699 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=396970 $D=8
XM753 24700 24701 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=431690 $D=8
XM754 24702 24703 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=432970 $D=8
XM755 24704 24705 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=467690 $D=8
XM756 23499 23500 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=468970 $D=8
XM757 VDD VSS VDD VDD pfet_03v3 L=2.505e-06 W=0.000166725 AD=0 AS=2.0381e-10 PD=0 PS=0.00079952 NRD=0 NRS=6.74977 m=1 nf=65 $X=146370 $Y=180915 $D=8
XM758 VDD 24106 23202 VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=156680 $Y=180895 $D=8
XM759 23209 24108 VDD VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=156680 $Y=213535 $D=8
XM760 VDD 24110 23210 VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=156680 $Y=216895 $D=8
XM761 23217 24112 VDD VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=156680 $Y=249535 $D=8
XM762 VDD 24114 23218 VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=156680 $Y=252895 $D=8
XM763 23225 24116 VDD VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=156680 $Y=285535 $D=8
XM764 VDD 24118 23226 VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=156680 $Y=288895 $D=8
XM765 23233 24120 VDD VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=156680 $Y=321535 $D=8
XM766 VDD 24122 23234 VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=156680 $Y=324895 $D=8
XM767 23241 24124 VDD VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=156680 $Y=357535 $D=8
XM768 VDD 24126 23242 VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=156680 $Y=360895 $D=8
XM769 23249 24128 VDD VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=156680 $Y=393535 $D=8
XM770 VDD 24130 23250 VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=156680 $Y=396895 $D=8
XM771 23257 24132 VDD VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=156680 $Y=429535 $D=8
XM772 VDD 24134 23258 VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=156680 $Y=432895 $D=8
XM773 23265 24136 VDD VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=156680 $Y=465535 $D=8
XM774 24043 1040 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=180895 $D=8
XM775 VDD 1044 24043 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=182015 $D=8
XM776 24043 1052 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=183135 $D=8
XM777 VDD 1045 24045 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=213535 $D=8
XM778 24045 1044 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=214655 $D=8
XM779 VDD 1040 24045 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=215775 $D=8
XM780 24047 1040 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=216895 $D=8
XM781 VDD 1043 24047 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=218015 $D=8
XM782 24047 1052 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=219135 $D=8
XM783 VDD 1045 24049 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=249535 $D=8
XM784 24049 1043 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=250655 $D=8
XM785 VDD 1040 24049 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=251775 $D=8
XM786 24051 1040 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=252895 $D=8
XM787 VDD 1042 24051 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=254015 $D=8
XM788 24051 1052 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=255135 $D=8
XM789 VDD 1045 24053 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=285535 $D=8
XM790 24053 1042 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=286655 $D=8
XM791 VDD 1040 24053 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=287775 $D=8
XM792 24055 1040 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=288895 $D=8
XM793 VDD 1041 24055 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=290015 $D=8
XM794 24055 1052 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=291135 $D=8
XM795 VDD 1045 24057 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=321535 $D=8
XM796 24057 1041 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=322655 $D=8
XM797 VDD 1040 24057 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=323775 $D=8
XM798 24059 1038 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=324895 $D=8
XM799 VDD 1044 24059 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=326015 $D=8
XM800 24059 1052 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=327135 $D=8
XM801 VDD 1045 24061 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=357535 $D=8
XM802 24061 1044 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=358655 $D=8
XM803 VDD 1038 24061 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=359775 $D=8
XM804 24063 1038 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=360895 $D=8
XM805 VDD 1043 24063 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=362015 $D=8
XM806 24063 1052 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=363135 $D=8
XM807 VDD 1045 24065 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=393535 $D=8
XM808 24065 1043 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=394655 $D=8
XM809 VDD 1038 24065 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=395775 $D=8
XM810 24067 1038 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=396895 $D=8
XM811 VDD 1042 24067 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=398015 $D=8
XM812 24067 1052 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=399135 $D=8
XM813 VDD 1045 24069 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=429535 $D=8
XM814 24069 1042 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=430655 $D=8
XM815 VDD 1038 24069 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=431775 $D=8
XM816 24071 1038 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=432895 $D=8
XM817 VDD 1041 24071 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=434015 $D=8
XM818 24071 1052 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=435135 $D=8
XM819 VDD 1045 24073 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=223995 $Y=465535 $D=8
XM820 24073 1041 VDD VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=223995 $Y=466655 $D=8
XM821 VDD 1038 24073 VDD pfet_03v3 L=2.8e-07 W=1.22e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=223995 $Y=467775 $D=8
XM822 24033 1 VDD VDD pfet_03v3 L=2.8e-07 W=1.06e-06 AD=5.985e-13 AS=1.3566e-12 PD=2.805e-06 PS=5.75e-06 NRD=0.115132 NRS=0.260965 m=1 nf=1 $X=233770 $Y=57780 $D=8
XM823 617 1000 VDD VDD pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=233770 $Y=63100 $D=8
XM824 1000 CLK 24033 VDD pfet_03v3 L=2.8e-07 W=1.06e-06 AD=1.3566e-12 AS=5.985e-13 PD=5.75e-06 PS=2.805e-06 NRD=0.260965 NRS=0.115132 m=1 nf=1 $X=234890 $Y=57780 $D=8
XM825 616 619 VDD VDD pfet_03v3 L=2.8e-07 W=5.29e-06 AD=2.9484e-12 AS=4.9896e-12 PD=1.238e-05 PS=2.444e-05 NRD=0.0917108 NRS=0.155203 m=1 nf=2 $X=242235 $Y=57810 $D=8
XM826 281 1006 VDD VDD pfet_03v3 L=4.65e-07 W=4.2e-07 AD=3.96e-13 AS=3.96e-13 PD=2.68e-06 PS=2.68e-06 NRD=0.488889 NRS=0.488889 m=1 nf=1 $X=243265 $Y=42525 $D=8
XM827 CEN 617 619 VDD pfet_03v3 L=2.8e-07 W=1.055e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=245925 $Y=59010 $D=8
XM828 618 1000 619 VDD pfet_03v3 L=2.8e-07 W=4.45e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=245925 $Y=64875 $D=8
XM829 317 281 VDD VDD pfet_03v3 L=2.8e-07 W=8.8e-07 AD=8.316e-13 AS=8.316e-13 PD=4.66e-06 PS=4.66e-06 NRD=0.232804 NRS=0.232804 m=1 nf=1 $X=246495 $Y=41535 $D=8
XM830 354 317 VDD VDD pfet_03v3 L=2.8e-07 W=3.515e-06 AD=1.9604e-12 AS=3.3176e-12 PD=8.58e-06 PS=1.684e-05 NRD=0.137931 NRS=0.233422 m=1 nf=2 $X=249065 $Y=39655 $D=8
XM831 250 468 VDD VDD pfet_03v3 L=2.8e-07 W=5.824e-5 AD=3.2448e-11 AS=3.69283e-11 PD=0.00013 PS=0.000130718 NRD=0.208333 NRS=0.237099 m=1 nf=10 $X=240535 $Y=94430 $D=8
XM832 445 354 VDD VDD pfet_03v3 L=2.8e-07 W=9.1e-06 AD=5.07e-12 AS=8.58e-12 PD=2.002e-05 PS=3.988e-05 NRD=0.0133333 NRS=0.0225641 m=1 nf=1 $X=256125 $Y=53590 $D=8
XM833 VDD CLK 445 VDD pfet_03v3 L=2.8e-07 W=9.1e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=257245 $Y=53590 $D=8
XM834 445 616 VDD VDD pfet_03v3 L=2.8e-07 W=9.1e-06 AD=8.58e-12 AS=5.07e-12 PD=3.988e-05 PS=2.002e-05 NRD=0.0225641 NRS=0.0133333 m=1 nf=1 $X=258365 $Y=53590 $D=8
XM835 VDD 495 468 VDD pfet_03v3 L=2.8e-07 W=1.058e-05 AD=5.8968e-12 AS=9.9792e-12 PD=2.32e-05 PS=4.624e-05 NRD=0.0114638 NRS=0.0194004 m=1 nf=1 $X=262120 $Y=50420 $D=8
XM836 468 445 VDD VDD pfet_03v3 L=2.8e-07 W=2.116e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.64e-05 PS=4.64e-05 NRD=0.0229277 NRS=0.0229277 m=1 nf=2 $X=263240 $Y=50420 $D=8
XM837 468 495 VDD VDD pfet_03v3 L=2.8e-07 W=1.058e-05 AD=9.9792e-12 AS=5.8968e-12 PD=4.624e-05 PS=2.32e-05 NRD=0.0194004 NRS=0.0114638 m=1 nf=1 $X=265480 $Y=50420 $D=8
XM838 VDD 24107 23266 VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=258945 $Y=180895 $D=8
XM839 23273 24109 VDD VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=258945 $Y=213535 $D=8
XM840 VDD 24111 23274 VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=258945 $Y=216895 $D=8
XM841 23281 24113 VDD VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=258945 $Y=249535 $D=8
XM842 VDD 24115 23282 VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=258945 $Y=252895 $D=8
XM843 23289 24117 VDD VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=258945 $Y=285535 $D=8
XM844 VDD 24119 23290 VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=258945 $Y=288895 $D=8
XM845 23297 24121 VDD VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=258945 $Y=321535 $D=8
XM846 VDD 24123 23298 VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=258945 $Y=324895 $D=8
XM847 23305 24125 VDD VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=258945 $Y=357535 $D=8
XM848 VDD 24127 23306 VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=258945 $Y=360895 $D=8
XM849 23313 24129 VDD VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=258945 $Y=393535 $D=8
XM850 VDD 24131 23314 VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=258945 $Y=396895 $D=8
XM851 23321 24133 VDD VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=258945 $Y=429535 $D=8
XM852 VDD 24135 23322 VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=258945 $Y=432895 $D=8
XM853 23329 24137 VDD VDD pfet_03v3 L=2.8e-07 W=1.4e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=258945 $Y=465535 $D=8
XM854 VDD 468 495 VDD pfet_03v3 L=2.8e-07 W=1.058e-05 AD=5.8968e-12 AS=9.9792e-12 PD=2.32e-05 PS=4.624e-05 NRD=0.0114638 NRS=0.0194004 m=1 nf=1 $X=268545 $Y=50420 $D=8
XM855 495 607 VDD VDD pfet_03v3 L=2.8e-07 W=2.116e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.64e-05 PS=4.64e-05 NRD=0.0229277 NRS=0.0229277 m=1 nf=2 $X=269665 $Y=50420 $D=8
XM856 495 468 VDD VDD pfet_03v3 L=2.8e-07 W=1.058e-05 AD=9.9792e-12 AS=5.8968e-12 PD=4.624e-05 PS=2.32e-05 NRD=0.0194004 NRS=0.0114638 m=1 nf=1 $X=271905 $Y=50420 $D=8
XM857 1 250 VDD VDD pfet_03v3 L=2.8e-07 W=1.7145e-04 AD=9.5524e-11 AS=1.02119e-10 PD=0.0003778 PS=0.000378518 NRD=0.28307 NRS=0.302613 m=1 nf=20 $X=253180 $Y=88540 $D=8
XM858 VDD VSS VDD VDD pfet_03v3 L=2.505e-06 W=0.000166725 AD=0 AS=2.0381e-10 PD=0 PS=0.00079952 NRD=0 NRS=6.74977 m=1 nf=65 $X=273750 $Y=180915 $D=8
XM859 VDD 23501 23502 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=179690 $D=8
XM860 VDD 24754 24755 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=180970 $D=8
XM861 VDD 24756 24757 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=215690 $D=8
XM862 VDD 24774 24775 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=216970 $D=8
XM863 VDD 24776 24777 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=251690 $D=8
XM864 VDD 24794 24795 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=252970 $D=8
XM865 VDD 24796 24797 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=287690 $D=8
XM866 VDD 24814 24815 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=288970 $D=8
XM867 VDD 24816 24817 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=323690 $D=8
XM868 VDD 24834 24835 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=324970 $D=8
XM869 VDD 24836 24837 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=359690 $D=8
XM870 VDD 24854 24855 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=360970 $D=8
XM871 VDD 24856 24857 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=395690 $D=8
XM872 VDD 24874 24875 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=396970 $D=8
XM873 VDD 24876 24877 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=431690 $D=8
XM874 VDD 24894 24895 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=432970 $D=8
XM875 VDD 24896 24897 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=467690 $D=8
XM876 VDD 23503 23504 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=468970 $D=8
XM877 23501 23502 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=179690 $D=8
XM878 24754 24755 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=180970 $D=8
XM879 24756 24757 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=215690 $D=8
XM880 24774 24775 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=216970 $D=8
XM881 24776 24777 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=251690 $D=8
XM882 24794 24795 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=252970 $D=8
XM883 24796 24797 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=287690 $D=8
XM884 24814 24815 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=288970 $D=8
XM885 24816 24817 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=323690 $D=8
XM886 24834 24835 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=324970 $D=8
XM887 24836 24837 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=359690 $D=8
XM888 24854 24855 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=360970 $D=8
XM889 24856 24857 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=395690 $D=8
XM890 24874 24875 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=396970 $D=8
XM891 24876 24877 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=431690 $D=8
XM892 24894 24895 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=432970 $D=8
XM893 24896 24897 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=467690 $D=8
XM894 23503 23504 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=468970 $D=8
XM895 VDD 23478 23480 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=179690 $D=8
XM896 VDD 24739 24738 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=180970 $D=8
XM897 VDD 24747 24746 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=215690 $D=8
XM898 VDD 24759 24758 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=216970 $D=8
XM899 VDD 24767 24766 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=251690 $D=8
XM900 VDD 24779 24778 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=252970 $D=8
XM901 VDD 24787 24786 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=287690 $D=8
XM902 VDD 24799 24798 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=288970 $D=8
XM903 VDD 24807 24806 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=323690 $D=8
XM904 VDD 24819 24818 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=324970 $D=8
XM905 VDD 24827 24826 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=359690 $D=8
XM906 VDD 24839 24838 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=360970 $D=8
XM907 VDD 24847 24846 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=395690 $D=8
XM908 VDD 24859 24858 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=396970 $D=8
XM909 VDD 24867 24866 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=431690 $D=8
XM910 VDD 24879 24878 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=432970 $D=8
XM911 VDD 24887 24886 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=467690 $D=8
XM912 VDD 23414 23416 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=468970 $D=8
XM913 23478 23480 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=179690 $D=8
XM914 24739 24738 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=180970 $D=8
XM915 24747 24746 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=215690 $D=8
XM916 24759 24758 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=216970 $D=8
XM917 24767 24766 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=251690 $D=8
XM918 24779 24778 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=252970 $D=8
XM919 24787 24786 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=287690 $D=8
XM920 24799 24798 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=288970 $D=8
XM921 24807 24806 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=323690 $D=8
XM922 24819 24818 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=324970 $D=8
XM923 24827 24826 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=359690 $D=8
XM924 24839 24838 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=360970 $D=8
XM925 24847 24846 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=395690 $D=8
XM926 24859 24858 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=396970 $D=8
XM927 24867 24866 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=431690 $D=8
XM928 24879 24878 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=432970 $D=8
XM929 24887 24886 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=467690 $D=8
XM930 23414 23416 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=468970 $D=8
XM931 23943 23200 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=311500 $Y=160970 $D=8
XM932 23944 23200 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=311500 $Y=164845 $D=8
XM933 24152 23886 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=311715 $Y=112830 $D=8
XM934 VDD 23474 23476 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=179690 $D=8
XM935 VDD 24741 24740 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=180970 $D=8
XM936 VDD 24749 24748 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=215690 $D=8
XM937 VDD 24761 24760 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=216970 $D=8
XM938 VDD 24769 24768 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=251690 $D=8
XM939 VDD 24781 24780 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=252970 $D=8
XM940 VDD 24789 24788 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=287690 $D=8
XM941 VDD 24801 24800 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=288970 $D=8
XM942 VDD 24809 24808 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=323690 $D=8
XM943 VDD 24821 24820 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=324970 $D=8
XM944 VDD 24829 24828 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=359690 $D=8
XM945 VDD 24841 24840 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=360970 $D=8
XM946 VDD 24849 24848 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=395690 $D=8
XM947 VDD 24861 24860 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=396970 $D=8
XM948 VDD 24869 24868 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=431690 $D=8
XM949 VDD 24881 24880 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=432970 $D=8
XM950 VDD 24889 24888 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=467690 $D=8
XM951 VDD 23410 23412 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=468970 $D=8
XM952 23474 23476 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=179690 $D=8
XM953 24741 24740 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=180970 $D=8
XM954 24749 24748 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=215690 $D=8
XM955 24761 24760 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=216970 $D=8
XM956 24769 24768 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=251690 $D=8
XM957 24781 24780 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=252970 $D=8
XM958 24789 24788 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=287690 $D=8
XM959 24801 24800 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=288970 $D=8
XM960 24809 24808 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=323690 $D=8
XM961 24821 24820 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=324970 $D=8
XM962 24829 24828 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=359690 $D=8
XM963 24841 24840 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=360970 $D=8
XM964 24849 24848 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=395690 $D=8
XM965 24861 24860 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=396970 $D=8
XM966 24869 24868 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=431690 $D=8
XM967 24881 24880 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=432970 $D=8
XM968 24889 24888 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=467690 $D=8
XM969 23410 23412 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=468970 $D=8
XM970 24153 23887 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=314245 $Y=112830 $D=8
XM971 23946 23200 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=314600 $Y=160970 $D=8
XM972 23945 23200 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=314600 $Y=164845 $D=8
XM973 VDD 23470 23472 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=179690 $D=8
XM974 VDD 24743 24742 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=180970 $D=8
XM975 VDD 24751 24750 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=215690 $D=8
XM976 VDD 24763 24762 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=216970 $D=8
XM977 VDD 24771 24770 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=251690 $D=8
XM978 VDD 24783 24782 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=252970 $D=8
XM979 VDD 24791 24790 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=287690 $D=8
XM980 VDD 24803 24802 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=288970 $D=8
XM981 VDD 24811 24810 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=323690 $D=8
XM982 VDD 24823 24822 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=324970 $D=8
XM983 VDD 24831 24830 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=359690 $D=8
XM984 VDD 24843 24842 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=360970 $D=8
XM985 VDD 24851 24850 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=395690 $D=8
XM986 VDD 24863 24862 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=396970 $D=8
XM987 VDD 24871 24870 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=431690 $D=8
XM988 VDD 24883 24882 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=432970 $D=8
XM989 VDD 24891 24890 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=467690 $D=8
XM990 VDD 23406 23408 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=468970 $D=8
XM991 23470 23472 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=179690 $D=8
XM992 24743 24742 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=180970 $D=8
XM993 24751 24750 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=215690 $D=8
XM994 24763 24762 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=216970 $D=8
XM995 24771 24770 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=251690 $D=8
XM996 24783 24782 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=252970 $D=8
XM997 24791 24790 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=287690 $D=8
XM998 24803 24802 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=288970 $D=8
XM999 24811 24810 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=323690 $D=8
XM1000 24823 24822 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=324970 $D=8
XM1001 24831 24830 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=359690 $D=8
XM1002 24843 24842 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=360970 $D=8
XM1003 24851 24850 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=395690 $D=8
XM1004 24863 24862 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=396970 $D=8
XM1005 24871 24870 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=431690 $D=8
XM1006 24883 24882 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=432970 $D=8
XM1007 24891 24890 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=467690 $D=8
XM1008 23406 23408 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=468970 $D=8
XM1009 23947 23200 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=317695 $Y=160970 $D=8
XM1010 23948 23200 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=317695 $Y=164845 $D=8
XM1011 24154 23888 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=317910 $Y=112830 $D=8
XM1012 VDD 23466 23468 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=179690 $D=8
XM1013 VDD 24745 24744 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=180970 $D=8
XM1014 VDD 24753 24752 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=215690 $D=8
XM1015 VDD 24765 24764 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=216970 $D=8
XM1016 VDD 24773 24772 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=251690 $D=8
XM1017 VDD 24785 24784 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=252970 $D=8
XM1018 VDD 24793 24792 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=287690 $D=8
XM1019 VDD 24805 24804 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=288970 $D=8
XM1020 VDD 24813 24812 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=323690 $D=8
XM1021 VDD 24825 24824 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=324970 $D=8
XM1022 VDD 24833 24832 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=359690 $D=8
XM1023 VDD 24845 24844 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=360970 $D=8
XM1024 VDD 24853 24852 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=395690 $D=8
XM1025 VDD 24865 24864 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=396970 $D=8
XM1026 VDD 24873 24872 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=431690 $D=8
XM1027 VDD 24885 24884 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=432970 $D=8
XM1028 VDD 24893 24892 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=467690 $D=8
XM1029 VDD 23402 23404 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=468970 $D=8
XM1030 23466 23468 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=179690 $D=8
XM1031 24745 24744 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=180970 $D=8
XM1032 24753 24752 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=215690 $D=8
XM1033 24765 24764 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=216970 $D=8
XM1034 24773 24772 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=251690 $D=8
XM1035 24785 24784 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=252970 $D=8
XM1036 24793 24792 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=287690 $D=8
XM1037 24805 24804 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=288970 $D=8
XM1038 24813 24812 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=323690 $D=8
XM1039 24825 24824 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=324970 $D=8
XM1040 24833 24832 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=359690 $D=8
XM1041 24845 24844 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=360970 $D=8
XM1042 24853 24852 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=395690 $D=8
XM1043 24865 24864 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=396970 $D=8
XM1044 24873 24872 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=431690 $D=8
XM1045 24885 24884 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=432970 $D=8
XM1046 24893 24892 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=467690 $D=8
XM1047 23402 23404 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=468970 $D=8
XM1048 24155 23889 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=320440 $Y=112830 $D=8
XM1049 23950 23200 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=320795 $Y=160970 $D=8
XM1050 23949 23200 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=320795 $Y=164845 $D=8
XM1051 VDD 23374 23376 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=179690 $D=8
XM1052 VDD 24455 24454 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=180970 $D=8
XM1053 VDD 24479 24478 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=323690 $D=8
XM1054 VDD 24503 24502 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=324970 $D=8
XM1055 VDD 24527 24526 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=467690 $D=8
XM1056 VDD 23430 23432 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=468970 $D=8
XM1057 23374 23376 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=179690 $D=8
XM1058 24455 24454 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=180970 $D=8
XM1059 24479 24478 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=323690 $D=8
XM1060 24503 24502 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=324970 $D=8
XM1061 24527 24526 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=467690 $D=8
XM1062 23430 23432 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=468970 $D=8
XM1063 23951 23200 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=323885 $Y=160970 $D=8
XM1064 23952 23200 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=323885 $Y=164845 $D=8
XM1065 24156 23890 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=324100 $Y=112830 $D=8
XM1066 VDD 23370 23372 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=179690 $D=8
XM1067 VDD 24457 24456 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=180970 $D=8
XM1068 VDD 24481 24480 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=323690 $D=8
XM1069 VDD 24505 24504 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=324970 $D=8
XM1070 VDD 24529 24528 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=467690 $D=8
XM1071 VDD 23426 23428 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=468970 $D=8
XM1072 23370 23372 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=179690 $D=8
XM1073 24457 24456 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=180970 $D=8
XM1074 24481 24480 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=323690 $D=8
XM1075 24505 24504 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=324970 $D=8
XM1076 24529 24528 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=467690 $D=8
XM1077 23426 23428 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=468970 $D=8
XM1078 24157 23891 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=326630 $Y=112830 $D=8
XM1079 23954 23200 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=326985 $Y=160970 $D=8
XM1080 23953 23200 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=326985 $Y=164845 $D=8
XM1081 VDD 23382 23384 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=179690 $D=8
XM1082 VDD 24459 24458 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=180970 $D=8
XM1083 VDD 24483 24482 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=323690 $D=8
XM1084 VDD 24507 24506 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=324970 $D=8
XM1085 VDD 24531 24530 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=467690 $D=8
XM1086 VDD 23422 23424 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=468970 $D=8
XM1087 23382 23384 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=179690 $D=8
XM1088 24459 24458 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=180970 $D=8
XM1089 24483 24482 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=323690 $D=8
XM1090 24507 24506 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=324970 $D=8
XM1091 24531 24530 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=467690 $D=8
XM1092 23422 23424 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=468970 $D=8
XM1093 23955 23200 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=330080 $Y=160970 $D=8
XM1094 23956 23200 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=330080 $Y=164845 $D=8
XM1095 24158 23892 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=330295 $Y=112830 $D=8
XM1096 VDD 23378 23380 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=179690 $D=8
XM1097 VDD 24461 24460 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=180970 $D=8
XM1098 VDD 24485 24484 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=323690 $D=8
XM1099 VDD 24509 24508 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=324970 $D=8
XM1100 VDD 24533 24532 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=467690 $D=8
XM1101 VDD 23418 23420 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=468970 $D=8
XM1102 23378 23380 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=179690 $D=8
XM1103 24461 24460 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=180970 $D=8
XM1104 24485 24484 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=323690 $D=8
XM1105 24509 24508 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=324970 $D=8
XM1106 24533 24532 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=467690 $D=8
XM1107 23418 23420 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=468970 $D=8
XM1108 24036 23893 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=332825 $Y=112830 $D=8
XM1109 1069 23200 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=333000 $Y=160970 $D=8
XM1110 1070 23200 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=333000 $Y=164845 $D=8
XM1111 1083 1081 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=336455 $Y=160970 $D=8
XM1112 1084 1081 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=336455 $Y=164845 $D=8
XM1113 VDD 23726 23728 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=179690 $D=8
XM1114 VDD 24476 24477 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=180970 $D=8
XM1115 VDD 24500 24501 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=323690 $D=8
XM1116 VDD 24524 24525 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=324970 $D=8
XM1117 VDD 24548 24549 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=467690 $D=8
XM1118 VDD 23758 23760 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=468970 $D=8
XM1119 24040 23886 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=336500 $Y=112830 $D=8
XM1120 23726 23728 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=179690 $D=8
XM1121 24476 24477 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=180970 $D=8
XM1122 24500 24501 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=323690 $D=8
XM1123 24524 24525 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=324970 $D=8
XM1124 24548 24549 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=467690 $D=8
XM1125 23758 23760 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=468970 $D=8
XM1126 24666 23887 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=339025 $Y=112830 $D=8
XM1127 24011 1081 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=339380 $Y=160970 $D=8
XM1128 24012 1081 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=339380 $Y=164845 $D=8
XM1129 VDD 23722 23724 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=179690 $D=8
XM1130 VDD 24474 24475 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=180970 $D=8
XM1131 VDD 24498 24499 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=323690 $D=8
XM1132 VDD 24522 24523 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=324970 $D=8
XM1133 VDD 24546 24547 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=467690 $D=8
XM1134 VDD 23754 23756 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=468970 $D=8
XM1135 23722 23724 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=179690 $D=8
XM1136 24474 24475 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=180970 $D=8
XM1137 24498 24499 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=323690 $D=8
XM1138 24522 24523 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=324970 $D=8
XM1139 24546 24547 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=467690 $D=8
XM1140 23754 23756 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=468970 $D=8
XM1141 24010 1081 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=342475 $Y=160970 $D=8
XM1142 24009 1081 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=342475 $Y=164845 $D=8
XM1143 VDD 23718 23720 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=179690 $D=8
XM1144 VDD 24472 24473 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=180970 $D=8
XM1145 VDD 24496 24497 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=323690 $D=8
XM1146 VDD 24520 24521 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=324970 $D=8
XM1147 VDD 24544 24545 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=467690 $D=8
XM1148 VDD 23750 23752 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=468970 $D=8
XM1149 24665 23888 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=342690 $Y=112830 $D=8
XM1150 23718 23720 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=179690 $D=8
XM1151 24472 24473 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=180970 $D=8
XM1152 24496 24497 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=323690 $D=8
XM1153 24520 24521 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=324970 $D=8
XM1154 24544 24545 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=467690 $D=8
XM1155 23750 23752 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=468970 $D=8
XM1156 24664 23889 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=345220 $Y=112830 $D=8
XM1157 24007 1081 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=345575 $Y=160970 $D=8
XM1158 24008 1081 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=345575 $Y=164845 $D=8
XM1159 VDD 23714 23716 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=179690 $D=8
XM1160 VDD 24470 24471 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=180970 $D=8
XM1161 VDD 24494 24495 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=323690 $D=8
XM1162 VDD 24518 24519 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=324970 $D=8
XM1163 VDD 24542 24543 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=467690 $D=8
XM1164 VDD 23746 23748 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=468970 $D=8
XM1165 23714 23716 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=179690 $D=8
XM1166 24470 24471 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=180970 $D=8
XM1167 24494 24495 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=323690 $D=8
XM1168 24518 24519 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=324970 $D=8
XM1169 24542 24543 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=467690 $D=8
XM1170 23746 23748 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=468970 $D=8
XM1171 VDD 23710 23712 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=179690 $D=8
XM1172 VDD 24468 24469 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=180970 $D=8
XM1173 VDD 24492 24493 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=323690 $D=8
XM1174 VDD 24516 24517 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=324970 $D=8
XM1175 VDD 24540 24541 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=467690 $D=8
XM1176 VDD 23742 23744 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=468970 $D=8
XM1177 24006 1081 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=348665 $Y=160970 $D=8
XM1178 24005 1081 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=348665 $Y=164845 $D=8
XM1179 24663 23890 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=348880 $Y=112830 $D=8
XM1180 23710 23712 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=179690 $D=8
XM1181 24468 24469 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=180970 $D=8
XM1182 24492 24493 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=323690 $D=8
XM1183 24516 24517 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=324970 $D=8
XM1184 24540 24541 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=467690 $D=8
XM1185 23742 23744 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=468970 $D=8
XM1186 24662 23891 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=351410 $Y=112830 $D=8
XM1187 VDD 23706 23708 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=179690 $D=8
XM1188 VDD 24466 24467 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=180970 $D=8
XM1189 VDD 24490 24491 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=323690 $D=8
XM1190 VDD 24514 24515 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=324970 $D=8
XM1191 VDD 24538 24539 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=467690 $D=8
XM1192 VDD 23738 23740 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=468970 $D=8
XM1193 24003 1081 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=351765 $Y=160970 $D=8
XM1194 24004 1081 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=351765 $Y=164845 $D=8
XM1195 23706 23708 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=179690 $D=8
XM1196 24466 24467 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=180970 $D=8
XM1197 24490 24491 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=323690 $D=8
XM1198 24514 24515 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=324970 $D=8
XM1199 24538 24539 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=467690 $D=8
XM1200 23738 23740 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=468970 $D=8
XM1201 VDD 23702 23704 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=179690 $D=8
XM1202 VDD 24464 24465 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=180970 $D=8
XM1203 VDD 24488 24489 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=323690 $D=8
XM1204 VDD 24512 24513 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=324970 $D=8
XM1205 VDD 24536 24537 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=467690 $D=8
XM1206 VDD 23734 23736 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=468970 $D=8
XM1207 24002 1081 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=354860 $Y=160970 $D=8
XM1208 24001 1081 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=354860 $Y=164845 $D=8
XM1209 24661 23892 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=355075 $Y=112830 $D=8
XM1210 23702 23704 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=179690 $D=8
XM1211 24464 24465 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=180970 $D=8
XM1212 24488 24489 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=323690 $D=8
XM1213 24512 24513 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=324970 $D=8
XM1214 24536 24537 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=467690 $D=8
XM1215 23734 23736 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=468970 $D=8
XM1216 VDD 23698 23700 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=179690 $D=8
XM1217 VDD 24462 24463 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=180970 $D=8
XM1218 VDD 24486 24487 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=323690 $D=8
XM1219 VDD 24510 24511 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=324970 $D=8
XM1220 VDD 24534 24535 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=467690 $D=8
XM1221 VDD 23730 23732 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=468970 $D=8
XM1222 24660 23893 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=357605 $Y=112830 $D=8
XM1223 23999 1081 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=357960 $Y=160970 $D=8
XM1224 24000 1081 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=357960 $Y=164845 $D=8
XM1225 23698 23700 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=179690 $D=8
XM1226 24462 24463 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=180970 $D=8
XM1227 24486 24487 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=323690 $D=8
XM1228 24510 24511 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=324970 $D=8
XM1229 24534 24535 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=467690 $D=8
XM1230 23730 23732 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=468970 $D=8
XM1231 VDD 23494 23496 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=179690 $D=8
XM1232 VDD 24231 24230 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=180970 $D=8
XM1233 VDD 24239 24238 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=323690 $D=8
XM1234 VDD 24247 24246 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=324970 $D=8
XM1235 VDD 24255 24254 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=467690 $D=8
XM1236 VDD 23790 23792 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=468970 $D=8
XM1237 23494 23496 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=179690 $D=8
XM1238 24231 24230 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=180970 $D=8
XM1239 24239 24238 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=323690 $D=8
XM1240 24247 24246 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=324970 $D=8
XM1241 24255 24254 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=467690 $D=8
XM1242 23790 23792 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=468970 $D=8
XM1243 23957 23201 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=365500 $Y=160970 $D=8
XM1244 23958 23201 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=365500 $Y=164845 $D=8
XM1245 24159 23886 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=365715 $Y=112830 $D=8
XM1246 VDD 23490 23492 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=179690 $D=8
XM1247 VDD 24233 24232 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=180970 $D=8
XM1248 VDD 24241 24240 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=323690 $D=8
XM1249 VDD 24249 24248 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=324970 $D=8
XM1250 VDD 24257 24256 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=467690 $D=8
XM1251 VDD 23786 23788 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=468970 $D=8
XM1252 23490 23492 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=179690 $D=8
XM1253 24233 24232 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=180970 $D=8
XM1254 24241 24240 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=323690 $D=8
XM1255 24249 24248 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=324970 $D=8
XM1256 24257 24256 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=467690 $D=8
XM1257 23786 23788 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=468970 $D=8
XM1258 24160 23887 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=368245 $Y=112830 $D=8
XM1259 23960 23201 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=368600 $Y=160970 $D=8
XM1260 23959 23201 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=368600 $Y=164845 $D=8
XM1261 VDD 23486 23488 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=179690 $D=8
XM1262 VDD 24235 24234 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=180970 $D=8
XM1263 VDD 24243 24242 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=323690 $D=8
XM1264 VDD 24251 24250 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=324970 $D=8
XM1265 VDD 24259 24258 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=467690 $D=8
XM1266 VDD 23782 23784 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=468970 $D=8
XM1267 23486 23488 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=179690 $D=8
XM1268 24235 24234 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=180970 $D=8
XM1269 24243 24242 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=323690 $D=8
XM1270 24251 24250 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=324970 $D=8
XM1271 24259 24258 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=467690 $D=8
XM1272 23782 23784 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=468970 $D=8
XM1273 23961 23201 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=371695 $Y=160970 $D=8
XM1274 23962 23201 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=371695 $Y=164845 $D=8
XM1275 24161 23888 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=371910 $Y=112830 $D=8
XM1276 VDD 23482 23484 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=179690 $D=8
XM1277 VDD 24237 24236 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=180970 $D=8
XM1278 VDD 24245 24244 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=323690 $D=8
XM1279 VDD 24253 24252 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=324970 $D=8
XM1280 VDD 24261 24260 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=467690 $D=8
XM1281 VDD 23778 23780 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=468970 $D=8
XM1282 23482 23484 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=179690 $D=8
XM1283 24237 24236 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=180970 $D=8
XM1284 24245 24244 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=323690 $D=8
XM1285 24253 24252 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=324970 $D=8
XM1286 24261 24260 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=467690 $D=8
XM1287 23778 23780 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=468970 $D=8
XM1288 24162 23889 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=374440 $Y=112830 $D=8
XM1289 23964 23201 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=374795 $Y=160970 $D=8
XM1290 23963 23201 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=374795 $Y=164845 $D=8
XM1291 VDD 23390 23392 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=179690 $D=8
XM1292 VDD 24551 24550 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=180970 $D=8
XM1293 VDD 24575 24574 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=323690 $D=8
XM1294 VDD 24599 24598 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=324970 $D=8
XM1295 VDD 24623 24622 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=467690 $D=8
XM1296 VDD 23774 23776 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=468970 $D=8
XM1297 23390 23392 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=179690 $D=8
XM1298 24551 24550 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=180970 $D=8
XM1299 24575 24574 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=323690 $D=8
XM1300 24599 24598 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=324970 $D=8
XM1301 24623 24622 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=467690 $D=8
XM1302 23774 23776 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=468970 $D=8
XM1303 23965 23201 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=377885 $Y=160970 $D=8
XM1304 23966 23201 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=377885 $Y=164845 $D=8
XM1305 24163 23890 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=378100 $Y=112830 $D=8
XM1306 VDD 23386 23388 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=179690 $D=8
XM1307 VDD 24553 24552 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=180970 $D=8
XM1308 VDD 24577 24576 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=323690 $D=8
XM1309 VDD 24601 24600 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=324970 $D=8
XM1310 VDD 24625 24624 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=467690 $D=8
XM1311 VDD 23770 23772 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=468970 $D=8
XM1312 23386 23388 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=179690 $D=8
XM1313 24553 24552 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=180970 $D=8
XM1314 24577 24576 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=323690 $D=8
XM1315 24601 24600 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=324970 $D=8
XM1316 24625 24624 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=467690 $D=8
XM1317 23770 23772 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=468970 $D=8
XM1318 24164 23891 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=380630 $Y=112830 $D=8
XM1319 23968 23201 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=380985 $Y=160970 $D=8
XM1320 23967 23201 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=380985 $Y=164845 $D=8
XM1321 VDD 23398 23400 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=179690 $D=8
XM1322 VDD 24555 24554 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=180970 $D=8
XM1323 VDD 24579 24578 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=323690 $D=8
XM1324 VDD 24603 24602 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=324970 $D=8
XM1325 VDD 24627 24626 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=467690 $D=8
XM1326 VDD 23766 23768 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=468970 $D=8
XM1327 23398 23400 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=179690 $D=8
XM1328 24555 24554 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=180970 $D=8
XM1329 24579 24578 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=323690 $D=8
XM1330 24603 24602 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=324970 $D=8
XM1331 24627 24626 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=467690 $D=8
XM1332 23766 23768 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=468970 $D=8
XM1333 23969 23201 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=384080 $Y=160970 $D=8
XM1334 23970 23201 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=384080 $Y=164845 $D=8
XM1335 24165 23892 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=384295 $Y=112830 $D=8
XM1336 VDD 23394 23396 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=179690 $D=8
XM1337 VDD 24557 24556 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=180970 $D=8
XM1338 VDD 24581 24580 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=323690 $D=8
XM1339 VDD 24605 24604 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=324970 $D=8
XM1340 VDD 24629 24628 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=467690 $D=8
XM1341 VDD 23762 23764 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=468970 $D=8
XM1342 23394 23396 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=179690 $D=8
XM1343 24557 24556 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=180970 $D=8
XM1344 24581 24580 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=323690 $D=8
XM1345 24605 24604 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=324970 $D=8
XM1346 24629 24628 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=467690 $D=8
XM1347 23762 23764 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=468970 $D=8
XM1348 24037 23893 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=386825 $Y=112830 $D=8
XM1349 1072 23201 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=387000 $Y=160970 $D=8
XM1350 1073 23201 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=387000 $Y=164845 $D=8
XM1351 1086 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=390455 $Y=160970 $D=8
XM1352 1087 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=390455 $Y=164845 $D=8
XM1353 VDD 23822 23824 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=179690 $D=8
XM1354 VDD 24572 24573 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=180970 $D=8
XM1355 VDD 24596 24597 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=323690 $D=8
XM1356 VDD 24620 24621 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=324970 $D=8
XM1357 VDD 24644 24645 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=467690 $D=8
XM1358 VDD 23854 23856 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=468970 $D=8
XM1359 24041 23886 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=390500 $Y=112830 $D=8
XM1360 23822 23824 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=179690 $D=8
XM1361 24572 24573 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=180970 $D=8
XM1362 24596 24597 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=323690 $D=8
XM1363 24620 24621 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=324970 $D=8
XM1364 24644 24645 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=467690 $D=8
XM1365 23854 23856 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=468970 $D=8
XM1366 24673 23887 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=393025 $Y=112830 $D=8
XM1367 24025 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=393380 $Y=160970 $D=8
XM1368 24026 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=393380 $Y=164845 $D=8
XM1369 VDD 23818 23820 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=179690 $D=8
XM1370 VDD 24570 24571 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=180970 $D=8
XM1371 VDD 24594 24595 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=323690 $D=8
XM1372 VDD 24618 24619 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=324970 $D=8
XM1373 VDD 24642 24643 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=467690 $D=8
XM1374 VDD 23850 23852 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=468970 $D=8
XM1375 23818 23820 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=179690 $D=8
XM1376 24570 24571 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=180970 $D=8
XM1377 24594 24595 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=323690 $D=8
XM1378 24618 24619 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=324970 $D=8
XM1379 24642 24643 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=467690 $D=8
XM1380 23850 23852 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=468970 $D=8
XM1381 24024 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=396475 $Y=160970 $D=8
XM1382 24023 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=396475 $Y=164845 $D=8
XM1383 VDD 23814 23816 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=179690 $D=8
XM1384 VDD 24568 24569 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=180970 $D=8
XM1385 VDD 24592 24593 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=323690 $D=8
XM1386 VDD 24616 24617 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=324970 $D=8
XM1387 VDD 24640 24641 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=467690 $D=8
XM1388 VDD 23846 23848 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=468970 $D=8
XM1389 24672 23888 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=396690 $Y=112830 $D=8
XM1390 23814 23816 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=179690 $D=8
XM1391 24568 24569 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=180970 $D=8
XM1392 24592 24593 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=323690 $D=8
XM1393 24616 24617 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=324970 $D=8
XM1394 24640 24641 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=467690 $D=8
XM1395 23846 23848 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=468970 $D=8
XM1396 24671 23889 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=399220 $Y=112830 $D=8
XM1397 24021 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=399575 $Y=160970 $D=8
XM1398 24022 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=399575 $Y=164845 $D=8
XM1399 VDD 23810 23812 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=179690 $D=8
XM1400 VDD 24566 24567 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=180970 $D=8
XM1401 VDD 24590 24591 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=323690 $D=8
XM1402 VDD 24614 24615 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=324970 $D=8
XM1403 VDD 24638 24639 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=467690 $D=8
XM1404 VDD 23842 23844 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=468970 $D=8
XM1405 23810 23812 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=179690 $D=8
XM1406 24566 24567 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=180970 $D=8
XM1407 24590 24591 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=323690 $D=8
XM1408 24614 24615 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=324970 $D=8
XM1409 24638 24639 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=467690 $D=8
XM1410 23842 23844 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=468970 $D=8
XM1411 VDD 23806 23808 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=179690 $D=8
XM1412 VDD 24564 24565 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=180970 $D=8
XM1413 VDD 24588 24589 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=323690 $D=8
XM1414 VDD 24612 24613 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=324970 $D=8
XM1415 VDD 24636 24637 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=467690 $D=8
XM1416 VDD 23838 23840 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=468970 $D=8
XM1417 24020 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=402665 $Y=160970 $D=8
XM1418 24019 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=402665 $Y=164845 $D=8
XM1419 24670 23890 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=402880 $Y=112830 $D=8
XM1420 23806 23808 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=179690 $D=8
XM1421 24564 24565 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=180970 $D=8
XM1422 24588 24589 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=323690 $D=8
XM1423 24612 24613 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=324970 $D=8
XM1424 24636 24637 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=467690 $D=8
XM1425 23838 23840 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=468970 $D=8
XM1426 24669 23891 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=405410 $Y=112830 $D=8
XM1427 VDD 23802 23804 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=179690 $D=8
XM1428 VDD 24562 24563 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=180970 $D=8
XM1429 VDD 24586 24587 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=323690 $D=8
XM1430 VDD 24610 24611 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=324970 $D=8
XM1431 VDD 24634 24635 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=467690 $D=8
XM1432 VDD 23834 23836 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=468970 $D=8
XM1433 24017 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=405765 $Y=160970 $D=8
XM1434 24018 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=405765 $Y=164845 $D=8
XM1435 23802 23804 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=179690 $D=8
XM1436 24562 24563 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=180970 $D=8
XM1437 24586 24587 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=323690 $D=8
XM1438 24610 24611 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=324970 $D=8
XM1439 24634 24635 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=467690 $D=8
XM1440 23834 23836 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=468970 $D=8
XM1441 VDD 23798 23800 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=179690 $D=8
XM1442 VDD 24560 24561 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=180970 $D=8
XM1443 VDD 24584 24585 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=323690 $D=8
XM1444 VDD 24608 24609 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=324970 $D=8
XM1445 VDD 24632 24633 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=467690 $D=8
XM1446 VDD 23830 23832 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=468970 $D=8
XM1447 24016 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=408860 $Y=160970 $D=8
XM1448 24015 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=408860 $Y=164845 $D=8
XM1449 24668 23892 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=409075 $Y=112830 $D=8
XM1450 23798 23800 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=179690 $D=8
XM1451 24560 24561 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=180970 $D=8
XM1452 24584 24585 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=323690 $D=8
XM1453 24608 24609 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=324970 $D=8
XM1454 24632 24633 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=467690 $D=8
XM1455 23830 23832 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=468970 $D=8
XM1456 VDD 23794 23796 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=179690 $D=8
XM1457 VDD 24558 24559 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=180970 $D=8
XM1458 VDD 24582 24583 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=323690 $D=8
XM1459 VDD 24606 24607 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=324970 $D=8
XM1460 VDD 24630 24631 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=467690 $D=8
XM1461 VDD 23826 23828 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=468970 $D=8
XM1462 24667 23893 VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=411605 $Y=112830 $D=8
XM1463 24013 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=411960 $Y=160970 $D=8
XM1464 24014 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=411960 $Y=164845 $D=8
XM1465 23794 23796 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=179690 $D=8
XM1466 24558 24559 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=180970 $D=8
XM1467 24582 24583 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=323690 $D=8
XM1468 24606 24607 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=324970 $D=8
XM1469 24630 24631 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=467690 $D=8
XM1470 23826 23828 VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=468970 $D=8
XM1471 VDD VSS VDD VDD pfet_03v3 L=1.74e-06 W=3.816e-05 AD=0 AS=6.1309e-11 PD=0 PS=0.000217698 NRD=0 NRS=11.8457 m=1 nf=36 $X=304360 $Y=171065 $D=8
XM1472 VDD VDD 23859 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=418720 $Y=467690 $D=8
XM1473 VDD VDD 23857 VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=418720 $Y=468970 $D=8
XM1474 614 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=6.35965e-12 PD=7.86e-06 PS=1.737e-05 NRD=0.152493 NRS=0.546921 m=1 nf=2 $X=418655 $Y=160970 $D=8
XM1475 615 1062 VDD VDD pfet_03v3 L=2.8e-07 W=3.18e-06 AD=1.7732e-12 AS=6.35965e-12 PD=7.86e-06 PS=1.737e-05 NRD=0.152493 NRS=0.546921 m=1 nf=2 $X=418655 $Y=164845 $D=8
XM1476 23860 VSS VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=419860 $Y=467690 $D=8
XM1477 23858 VSS VDD VDD pfet_03v3 L=2.8e-07 W=2.8e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=419860 $Y=468970 $D=8
XM1478 606 614 VDD VDD pfet_03v3 L=2.8e-07 W=3.275e-06 AD=1.8252e-12 AS=3.0888e-12 PD=8.06e-06 PS=1.58e-05 NRD=0.148148 NRS=0.250712 m=1 nf=2 $X=418770 $Y=97440 $D=8
XM1479 607 606 VDD VDD pfet_03v3 L=2.8e-07 W=9.93e-06 AD=5.5328e-12 AS=9.3632e-12 PD=2.232e-05 PS=4.432e-05 NRD=0.0488722 NRS=0.0827068 m=1 nf=2 $X=418790 $Y=67070 $D=8
XM1480 613 VDD VDD VDD pfet_03v3 L=2.8e-07 W=1.385e-06 AD=9.801e-13 AS=2.33887e-12 PD=4.29e-06 PS=9.09e-06 NRD=0.444444 NRS=1.06061 m=1 nf=2 $X=418870 $Y=112830 $D=8
X1488 614 614 613 VDD pfet_03v3_I13 $T=419815 124190 0 180 $X=418175 $Y=116760
X1489 615 615 613 VDD pfet_03v3_I13 $T=419815 151940 0 180 $X=418175 $Y=144510
X1490 615 614 1062 VDD pfet_03v3_I13 $T=419825 159875 0 180 $X=418185 $Y=152445
X1491 614 614 VDD VSS nfet_03v3_I02 $T=419815 133465 0 180 $X=418535 $Y=126035
X1492 615 615 VDD VSS nfet_03v3_I02 $T=419815 143485 0 180 $X=418535 $Y=136055
X1498 VDD 618 616 pmos_1p2$$46273580 $T=242390 65835 1 0 $X=240960 $Y=64015
X1499 VSS 617 1000 VSS nmos_1p2$$46563372 $T=233925 66830 0 0 $X=232780 $Y=66145
X1500 618 VSS 616 VSS nmos_1p2$$46563372 $T=243510 68190 1 0 $X=242365 $Y=66555
X1501 619 618 617 VSS nmos_1p2$$46563372 $T=246080 68190 1 0 $X=244935 $Y=66555
X1503 1063 VSS Q[0] D[0] 23198 1 VDD 1064 1065 WEN[0] 23915 23916 23917 23918 23919 23920 23921 23922 23923 23924
+ 23925 23926 23927 23928 24034 1053 23885 23884 23883 23882 23881 23880 23879 23878 23877 24138 24139 24140 24141 24142
+ 24143 24144
+ saout_m2 $T=9775 25090 0 0 $X=8430 $Y=7315
X1504 1032 VSS Q[2] D[2] 23199 1 VDD 1066 1067 WEN[2] 23929 23930 23931 23932 23933 23934 23935 23936 23937 23938
+ 23939 23940 23941 23942 24035 1053 23885 23884 23883 23882 23881 23880 23879 23878 23877 24145 24146 24147 24148 24149
+ 24150 24151
+ saout_m2 $T=63775 25090 0 0 $X=62430 $Y=7315
X1505 1068 VSS Q[4] D[4] 23200 1 VDD 1069 1070 WEN[4] 23943 23944 23945 23946 23947 23948 23949 23950 23951 23952
+ 23953 23954 23955 23956 24036 1053 23886 23887 23888 23889 23890 23891 23892 23893 23877 24152 24153 24154 24155 24156
+ 24157 24158
+ saout_m2 $T=307655 25090 0 0 $X=306310 $Y=7315
X1506 1071 VSS Q[6] D[6] 23201 1 VDD 1072 1073 WEN[6] 23957 23958 23959 23960 23961 23962 23963 23964 23965 23966
+ 23967 23968 23969 23970 24037 1053 23886 23887 23888 23889 23890 23891 23892 23893 23877 24159 24160 24161 24162 24163
+ 24164 24165
+ saout_m2 $T=361655 25090 0 0 $X=360310 $Y=7315
X1507 VSS VSS 23337 23338 23339 23340 23341 23342 23343 23344 ICV_7 $T=27210 176130 1 180 $X=23870 $Y=175790
X1508 VSS VSS 23345 23346 23347 23348 23349 23350 23351 23352 ICV_7 $T=33210 176130 1 180 $X=29870 $Y=175790
X1509 VSS VSS 23353 23354 23355 23356 23357 23358 23359 23360 ICV_7 $T=81210 176130 1 180 $X=77870 $Y=175790
X1510 VSS VSS 23361 23362 23363 23364 23365 23366 23367 23368 ICV_7 $T=87210 176130 1 180 $X=83870 $Y=175790
X1511 VSS VSS 23369 23370 23371 23372 23373 23374 23375 23376 ICV_7 $T=325090 176130 1 180 $X=321750 $Y=175790
X1512 VSS VSS 23377 23378 23379 23380 23381 23382 23383 23384 ICV_7 $T=331090 176130 1 180 $X=327750 $Y=175790
X1513 VSS VSS 23385 23386 23387 23388 23389 23390 23391 23392 ICV_7 $T=379090 176130 1 180 $X=375750 $Y=175790
X1514 VSS VSS 23393 23394 23395 23396 23397 23398 23399 23400 ICV_7 $T=385090 176130 1 180 $X=381750 $Y=175790
X1515 VSS 1002 23401 23402 23403 23404 23405 23406 23407 23408 23409 23410 23411 23412 23413 23414 23415 23416 ICV_8 $T=313090 473130 0 180 $X=309750 $Y=468290
X1516 VSS 1002 23417 23418 23419 23420 23421 23422 23423 23424 23425 23426 23427 23428 23429 23430 23431 23432 ICV_8 $T=325090 473130 0 180 $X=321750 $Y=468290
X1520 VSS VSS 23433 23434 23435 23436 23437 23438 23439 23440 23441 23442 23443 23444 23445 23446 23447 23448 ICV_9 $T=12210 176130 1 180 $X=8870 $Y=175790
X1521 VSS VSS 23449 23450 23451 23452 23453 23454 23455 23456 23457 23458 23459 23460 23461 23462 23463 23464 ICV_9 $T=66210 176130 1 180 $X=62870 $Y=175790
X1522 VSS VSS 23465 23466 23467 23468 23469 23470 23471 23472 23473 23474 23475 23476 23477 23478 23479 23480 ICV_9 $T=310090 176130 1 180 $X=306750 $Y=175790
X1523 VSS VSS 23481 23482 23483 23484 23485 23486 23487 23488 23489 23490 23491 23492 23493 23494 23495 23496 ICV_9 $T=364090 176130 1 180 $X=360750 $Y=175790
X1528 VDD VSS 23202 23203 23204 23205 23206 23207 23208 23209 23210 23211 23212 23213 23214 23215 23216 23217 23218 23219
+ 23220 23221 23222 23223 23224 23225 23226 23227 23228 23229 23230 23231 23232 23233 23922 23921 23920 23919 23918 23917
+ 23916 23915 24166 24167 24168 24169 24170 24171 24172 24173 24174 24175 24176 24177 24178 24179 24180 24181
+ ICV_27 $T=12210 185130 1 180 $X=8870 $Y=180290
X1529 VDD VSS 23234 23235 23236 23237 23238 23239 23240 23241 23242 23243 23244 23245 23246 23247 23248 23249 23250 23251
+ 23252 23253 23254 23255 23256 23257 23258 23259 23260 23261 23262 23263 23264 23265 23922 23921 23920 23919 23918 23917
+ 23916 23915 24182 24183 24184 24185 24186 24187 24188 24189 24190 24191 24192 24193 24194 24195 24196 24197
+ ICV_27 $T=12210 329130 1 180 $X=8870 $Y=324290
X1530 VDD VSS 23202 23203 23204 23205 23206 23207 23208 23209 23210 23211 23212 23213 23214 23215 23216 23217 23218 23219
+ 23220 23221 23222 23223 23224 23225 23226 23227 23228 23229 23230 23231 23232 23233 23936 23935 23934 23933 23932 23931
+ 23930 23929 24198 24199 24200 24201 24202 24203 24204 24205 24206 24207 24208 24209 24210 24211 24212 24213
+ ICV_27 $T=66210 185130 1 180 $X=62870 $Y=180290
X1531 VDD VSS 23234 23235 23236 23237 23238 23239 23240 23241 23242 23243 23244 23245 23246 23247 23248 23249 23250 23251
+ 23252 23253 23254 23255 23256 23257 23258 23259 23260 23261 23262 23263 23264 23265 23936 23935 23934 23933 23932 23931
+ 23930 23929 24214 24215 24216 24217 24218 24219 24220 24221 24222 24223 24224 24225 24226 24227 24228 24229
+ ICV_27 $T=66210 329130 1 180 $X=62870 $Y=324290
X1532 VDD VSS 23266 23267 23268 23269 23270 23271 23272 23273 23274 23275 23276 23277 23278 23279 23280 23281 23282 23283
+ 23284 23285 23286 23287 23288 23289 23290 23291 23292 23293 23294 23295 23296 23297 23964 23963 23962 23961 23960 23959
+ 23958 23957 24230 24231 24232 24233 24234 24235 24236 24237 24238 24239 24240 24241 24242 24243 24244 24245
+ ICV_27 $T=364090 185130 1 180 $X=360750 $Y=180290
X1533 VDD VSS 23298 23299 23300 23301 23302 23303 23304 23305 23306 23307 23308 23309 23310 23311 23312 23313 23314 23315
+ 23316 23317 23318 23319 23320 23321 23322 23323 23324 23325 23326 23327 23328 23329 23964 23963 23962 23961 23960 23959
+ 23958 23957 24246 24247 24248 24249 24250 24251 24252 24253 24254 24255 24256 24257 24258 24259 24260 24261
+ ICV_27 $T=364090 329130 1 180 $X=360750 $Y=324290
X1534 VSS VSS 23505 23506 23507 23508 23509 23510 23511 23512 23513 23514 23515 23516 23517 23518 23519 23520 23521 23522
+ 23523 23524 23525 23526 23527 23528 23529 23530 23531 23532 23533 23534 23535 23536
+ ICV_10 $T=12210 473130 0 180 $X=8870 $Y=468290
X1535 VSS VSS 23537 23538 23539 23540 23541 23542 23543 23544 23545 23546 23547 23548 23549 23550 23551 23552 23553 23554
+ 23555 23556 23557 23558 23559 23560 23561 23562 23563 23564 23565 23566 23567 23568
+ ICV_10 $T=39210 176130 1 180 $X=35870 $Y=175790
X1536 VSS VSS 23569 23570 23571 23572 23573 23574 23575 23576 23577 23578 23579 23580 23581 23582 23583 23584 23585 23586
+ 23587 23588 23589 23590 23591 23592 23593 23594 23595 23596 23597 23598 23599 23600
+ ICV_10 $T=39210 473130 0 180 $X=35870 $Y=468290
X1537 VSS VSS 23601 23602 23603 23604 23605 23606 23607 23608 23609 23610 23611 23612 23613 23614 23615 23616 23617 23618
+ 23619 23620 23621 23622 23623 23624 23625 23626 23627 23628 23629 23630 23631 23632
+ ICV_10 $T=66210 473130 0 180 $X=62870 $Y=468290
X1538 VSS VSS 23633 23634 23635 23636 23637 23638 23639 23640 23641 23642 23643 23644 23645 23646 23647 23648 23649 23650
+ 23651 23652 23653 23654 23655 23656 23657 23658 23659 23660 23661 23662 23663 23664
+ ICV_10 $T=93210 176130 1 180 $X=89870 $Y=175790
X1539 VSS VSS 23665 23666 23667 23668 23669 23670 23671 23672 23673 23674 23675 23676 23677 23678 23679 23680 23681 23682
+ 23683 23684 23685 23686 23687 23688 23689 23690 23691 23692 23693 23694 23695 23696
+ ICV_10 $T=93210 473130 0 180 $X=89870 $Y=468290
X1540 VSS VSS 23697 23698 23699 23700 23701 23702 23703 23704 23705 23706 23707 23708 23709 23710 23711 23712 23713 23714
+ 23715 23716 23717 23718 23719 23720 23721 23722 23723 23724 23725 23726 23727 23728
+ ICV_10 $T=337090 176130 1 180 $X=333750 $Y=175790
X1541 VSS 1002 23729 23730 23731 23732 23733 23734 23735 23736 23737 23738 23739 23740 23741 23742 23743 23744 23745 23746
+ 23747 23748 23749 23750 23751 23752 23753 23754 23755 23756 23757 23758 23759 23760
+ ICV_10 $T=337090 473130 0 180 $X=333750 $Y=468290
X1542 VSS 1002 23761 23762 23763 23764 23765 23766 23767 23768 23769 23770 23771 23772 23773 23774 23775 23776 23777 23778
+ 23779 23780 23781 23782 23783 23784 23785 23786 23787 23788 23789 23790 23791 23792
+ ICV_10 $T=364090 473130 0 180 $X=360750 $Y=468290
X1543 VSS VSS 23793 23794 23795 23796 23797 23798 23799 23800 23801 23802 23803 23804 23805 23806 23807 23808 23809 23810
+ 23811 23812 23813 23814 23815 23816 23817 23818 23819 23820 23821 23822 23823 23824
+ ICV_10 $T=391090 176130 1 180 $X=387750 $Y=175790
X1544 VSS 1002 23825 23826 23827 23828 23829 23830 23831 23832 23833 23834 23835 23836 23837 23838 23839 23840 23841 23842
+ 23843 23844 23845 23846 23847 23848 23849 23850 23851 23852 23853 23854 23855 23856
+ ICV_10 $T=391090 473130 0 180 $X=387750 $Y=468290
X1568 VDD VSS 23202 23203 23204 23205 23206 23207 23208 23209 23210 23211 23212 23213 23214 23215 23216 23217 23218 23219
+ 23220 23221 23222 23223 23224 23225 23226 23227 23228 23229 23230 23231 23232 23233 23923 23924 23925 23926 23927 23928
+ 1065 1064 1076 1077 23984 23983 23982 23981 23980 23979 23978 23977 23976 23975 23974 23973 23972 23971 24262 24263
+ 24264 24265 24266 24267 24268 24269 24270 24271 24272 24273 24274 24275 24276 24277 24278 24279 24280 24281 24282 24283
+ 24284 24285 24286 24287 24288 24289 24290 24291 24292 24293 24294 24295 24296 24297 24298 24299 24300 24301 24302 24303
+ 24304 24305 24306 24307 24308 24309
+ ICV_24 $T=24210 180630 0 0 $X=23870 $Y=180290
X1569 VDD VSS 23234 23235 23236 23237 23238 23239 23240 23241 23242 23243 23244 23245 23246 23247 23248 23249 23250 23251
+ 23252 23253 23254 23255 23256 23257 23258 23259 23260 23261 23262 23263 23264 23265 23923 23924 23925 23926 23927 23928
+ 1065 1064 1076 1077 23984 23983 23982 23981 23980 23979 23978 23977 23976 23975 23974 23973 23972 23971 24310 24311
+ 24312 24313 24314 24315 24316 24317 24318 24319 24320 24321 24322 24323 24324 24325 24326 24327 24328 24329 24330 24331
+ 24332 24333 24334 24335 24336 24337 24338 24339 24340 24341 24342 24343 24344 24345 24346 24347 24348 24349 24350 24351
+ 24352 24353 24354 24355 24356 24357
+ ICV_24 $T=24210 324630 0 0 $X=23870 $Y=324290
X1570 VDD VSS 23202 23203 23204 23205 23206 23207 23208 23209 23210 23211 23212 23213 23214 23215 23216 23217 23218 23219
+ 23220 23221 23222 23223 23224 23225 23226 23227 23228 23229 23230 23231 23232 23233 23937 23938 23939 23940 23941 23942
+ 1067 1066 1079 1080 23998 23997 23996 23995 23994 23993 23992 23991 23990 23989 23988 23987 23986 23985 24358 24359
+ 24360 24361 24362 24363 24364 24365 24366 24367 24368 24369 24370 24371 24372 24373 24374 24375 24376 24377 24378 24379
+ 24380 24381 24382 24383 24384 24385 24386 24387 24388 24389 24390 24391 24392 24393 24394 24395 24396 24397 24398 24399
+ 24400 24401 24402 24403 24404 24405
+ ICV_24 $T=78210 180630 0 0 $X=77870 $Y=180290
X1571 VDD VSS 23234 23235 23236 23237 23238 23239 23240 23241 23242 23243 23244 23245 23246 23247 23248 23249 23250 23251
+ 23252 23253 23254 23255 23256 23257 23258 23259 23260 23261 23262 23263 23264 23265 23937 23938 23939 23940 23941 23942
+ 1067 1066 1079 1080 23998 23997 23996 23995 23994 23993 23992 23991 23990 23989 23988 23987 23986 23985 24406 24407
+ 24408 24409 24410 24411 24412 24413 24414 24415 24416 24417 24418 24419 24420 24421 24422 24423 24424 24425 24426 24427
+ 24428 24429 24430 24431 24432 24433 24434 24435 24436 24437 24438 24439 24440 24441 24442 24443 24444 24445 24446 24447
+ 24448 24449 24450 24451 24452 24453
+ ICV_24 $T=78210 324630 0 0 $X=77870 $Y=324290
X1572 VDD VSS 23266 23267 23268 23269 23270 23271 23272 23273 23274 23275 23276 23277 23278 23279 23280 23281 23282 23283
+ 23284 23285 23286 23287 23288 23289 23290 23291 23292 23293 23294 23295 23296 23297 23951 23952 23953 23954 23955 23956
+ 1070 1069 1083 1084 24012 24011 24010 24009 24008 24007 24006 24005 24004 24003 24002 24001 24000 23999 24454 24455
+ 24456 24457 24458 24459 24460 24461 24462 24463 24464 24465 24466 24467 24468 24469 24470 24471 24472 24473 24474 24475
+ 24476 24477 24478 24479 24480 24481 24482 24483 24484 24485 24486 24487 24488 24489 24490 24491 24492 24493 24494 24495
+ 24496 24497 24498 24499 24500 24501
+ ICV_24 $T=322090 180630 0 0 $X=321750 $Y=180290
X1573 VDD VSS 23298 23299 23300 23301 23302 23303 23304 23305 23306 23307 23308 23309 23310 23311 23312 23313 23314 23315
+ 23316 23317 23318 23319 23320 23321 23322 23323 23324 23325 23326 23327 23328 23329 23951 23952 23953 23954 23955 23956
+ 1070 1069 1083 1084 24012 24011 24010 24009 24008 24007 24006 24005 24004 24003 24002 24001 24000 23999 24502 24503
+ 24504 24505 24506 24507 24508 24509 24510 24511 24512 24513 24514 24515 24516 24517 24518 24519 24520 24521 24522 24523
+ 24524 24525 24526 24527 24528 24529 24530 24531 24532 24533 24534 24535 24536 24537 24538 24539 24540 24541 24542 24543
+ 24544 24545 24546 24547 24548 24549
+ ICV_24 $T=322090 324630 0 0 $X=321750 $Y=324290
X1574 VDD VSS 23266 23267 23268 23269 23270 23271 23272 23273 23274 23275 23276 23277 23278 23279 23280 23281 23282 23283
+ 23284 23285 23286 23287 23288 23289 23290 23291 23292 23293 23294 23295 23296 23297 23965 23966 23967 23968 23969 23970
+ 1073 1072 1086 1087 24026 24025 24024 24023 24022 24021 24020 24019 24018 24017 24016 24015 24014 24013 24550 24551
+ 24552 24553 24554 24555 24556 24557 24558 24559 24560 24561 24562 24563 24564 24565 24566 24567 24568 24569 24570 24571
+ 24572 24573 24574 24575 24576 24577 24578 24579 24580 24581 24582 24583 24584 24585 24586 24587 24588 24589 24590 24591
+ 24592 24593 24594 24595 24596 24597
+ ICV_24 $T=376090 180630 0 0 $X=375750 $Y=180290
X1575 VDD VSS 23298 23299 23300 23301 23302 23303 23304 23305 23306 23307 23308 23309 23310 23311 23312 23313 23314 23315
+ 23316 23317 23318 23319 23320 23321 23322 23323 23324 23325 23326 23327 23328 23329 23965 23966 23967 23968 23969 23970
+ 1073 1072 1086 1087 24026 24025 24024 24023 24022 24021 24020 24019 24018 24017 24016 24015 24014 24013 24598 24599
+ 24600 24601 24602 24603 24604 24605 24606 24607 24608 24609 24610 24611 24612 24613 24614 24615 24616 24617 24618 24619
+ 24620 24621 24622 24623 24624 24625 24626 24627 24628 24629 24630 24631 24632 24633 24634 24635 24636 24637 24638 24639
+ 24640 24641 24642 24643 24644 24645
+ ICV_24 $T=376090 324630 0 0 $X=375750 $Y=324290
X1576 1075 VSS Q[1] 1074 D[1] 1 VDD 1076 1077 WEN[1] 23971 23972 23973 23974 23975 23976 23977 23978 23979 23980
+ 23981 23982 23983 23984 24038 1053 23878 23879 23880 23881 23882 23883 23884 23885 23877 24646 24647 24648 24649 24650
+ 24651 24652
+ saout_R_m2 $T=65645 25125 1 180 $X=27480 $Y=6815
X1577 1033 VSS Q[3] 1078 D[3] 1 VDD 1079 1080 WEN[3] 23985 23986 23987 23988 23989 23990 23991 23992 23993 23994
+ 23995 23996 23997 23998 24039 1053 23878 23879 23880 23881 23882 23883 23884 23885 23877 24653 24654 24655 24656 24657
+ 24658 24659
+ saout_R_m2 $T=119645 25125 1 180 $X=81480 $Y=6815
X1578 1082 VSS Q[5] 1081 D[5] 1 VDD 1083 1084 WEN[5] 23999 24000 24001 24002 24003 24004 24005 24006 24007 24008
+ 24009 24010 24011 24012 24040 1053 23893 23892 23891 23890 23889 23888 23887 23886 23877 24660 24661 24662 24663 24664
+ 24665 24666
+ saout_R_m2 $T=363525 25125 1 180 $X=325360 $Y=6815
X1579 1085 VSS Q[7] 1062 D[7] 1 VDD 1086 1087 WEN[7] 24013 24014 24015 24016 24017 24018 24019 24020 24021 24022
+ 24023 24024 24025 24026 24041 1053 23893 23892 23891 23890 23889 23888 23887 23886 23877 24667 24668 24669 24670 24671
+ 24672 24673
+ saout_R_m2 $T=417525 25125 1 180 $X=379360 $Y=6815
X1581 VDD VSS 702 703 24674 24675 24676 24677 ICV_41 $T=117210 185130 0 0 $X=116870 $Y=180290
X1582 VDD VSS 702 703 24678 24679 24680 24681 ICV_41 $T=117210 221130 0 0 $X=116870 $Y=216290
X1583 VDD VSS 702 703 24682 24683 24684 24685 ICV_41 $T=117210 257130 0 0 $X=116870 $Y=252290
X1584 VDD VSS 702 703 24686 24687 24688 24689 ICV_41 $T=117210 293130 0 0 $X=116870 $Y=288290
X1585 VDD VSS 702 703 24690 24691 24692 24693 ICV_41 $T=117210 329130 0 0 $X=116870 $Y=324290
X1586 VDD VSS 702 703 24694 24695 24696 24697 ICV_41 $T=117210 365130 0 0 $X=116870 $Y=360290
X1587 VDD VSS 702 703 24698 24699 24700 24701 ICV_41 $T=117210 401130 0 0 $X=116870 $Y=396290
X1588 VDD VSS 702 703 24702 24703 24704 24705 ICV_41 $T=117210 437130 0 0 $X=116870 $Y=432290
X1589 VSS VDD 1040 1044 1046 1047 1048 1049 1050 1051 23203 23204 23205 23206 23207 23208 23267 23268 23269 23270
+ 23271 23272 1 24042 24043 24044 24045 24106 24107 24108 24109
+ ICV_37 $T=154400 190385 1 270 $X=126565 $Y=179495
X1590 VSS VDD 1040 1043 1046 1047 1048 1049 1050 1051 23211 23212 23213 23214 23215 23216 23275 23276 23277 23278
+ 23279 23280 1 24046 24047 24048 24049 24110 24111 24112 24113
+ ICV_37 $T=154400 226385 1 270 $X=126565 $Y=215495
X1591 VSS VDD 1040 1042 1046 1047 1048 1049 1050 1051 23219 23220 23221 23222 23223 23224 23283 23284 23285 23286
+ 23287 23288 1 24050 24051 24052 24053 24114 24115 24116 24117
+ ICV_37 $T=154400 262385 1 270 $X=126565 $Y=251495
X1592 VSS VDD 1040 1041 1046 1047 1048 1049 1050 1051 23227 23228 23229 23230 23231 23232 23291 23292 23293 23294
+ 23295 23296 1 24054 24055 24056 24057 24118 24119 24120 24121
+ ICV_37 $T=154400 298385 1 270 $X=126565 $Y=287495
X1593 VSS VDD 1038 1044 1046 1047 1048 1049 1050 1051 23235 23236 23237 23238 23239 23240 23299 23300 23301 23302
+ 23303 23304 1 24058 24059 24060 24061 24122 24123 24124 24125
+ ICV_37 $T=154400 334385 1 270 $X=126565 $Y=323495
X1594 VSS VDD 1038 1043 1046 1047 1048 1049 1050 1051 23243 23244 23245 23246 23247 23248 23307 23308 23309 23310
+ 23311 23312 1 24062 24063 24064 24065 24126 24127 24128 24129
+ ICV_37 $T=154400 370385 1 270 $X=126565 $Y=359495
X1595 VSS VDD 1038 1042 1046 1047 1048 1049 1050 1051 23251 23252 23253 23254 23255 23256 23315 23316 23317 23318
+ 23319 23320 1 24066 24067 24068 24069 24130 24131 24132 24133
+ ICV_37 $T=154400 406385 1 270 $X=126565 $Y=395495
X1596 VSS VDD 1038 1041 1046 1047 1048 1049 1050 1051 23259 23260 23261 23262 23263 23264 23323 23324 23325 23326
+ 23327 23328 1 24070 24071 24072 24073 24134 24135 24136 24137
+ ICV_37 $T=154400 442385 1 270 $X=126565 $Y=431495
X1600 VSS VDD 1 CLK VSS A[8] 23902 23903 1038 1040 xpredec0 $T=146075 111460 0 0 $X=144630 $Y=111455
X1601 VSS VDD 1 CLK A[7] A[6] 1041 1042 1043 1044 xpredec0 $T=182970 111460 0 0 $X=181525 $Y=111455
X1606 VSS VDD 1 CLK 23884 23885 23878 23879 23880 23881 23882 23883 23893 23892 23891 23890 23889 23888 23887 23886
+ A[2] A[1] A[0]
+ ypredec1 $T=145470 26355 0 0 $X=146365 $Y=26735
X1609 1001 VSS 1003 nfet_03v3_I20 $T=175115 470995 0 90 $X=164385 $Y=470315
X1610 1002 VSS 1004 nfet_03v3_I20 $T=260115 470995 0 90 $X=249385 $Y=470315
X1614 VDD 1001 1003 pmos_1p2_02_R90 $T=189610 471150 0 90 $X=176320 $Y=469670
X1615 VDD 1002 1004 pmos_1p2_02_R90 $T=248135 471150 0 90 $X=234845 $Y=469670
X1616 1003 VDD 2 VDD pfet_03v3_I14 $T=198405 470995 0 90 $X=191195 $Y=469955
X1617 1 2 VSS VDD pfet_03v3_I14 $T=219905 470995 0 90 $X=212695 $Y=469955
X1618 1004 VDD 2 VDD pfet_03v3_I14 $T=233255 470995 0 90 $X=226045 $Y=469955
X1619 1003 VSS 2 nfet_03v3_I11 $T=202950 470995 0 90 $X=199690 $Y=470315
X1620 1004 VSS 2 nfet_03v3_I11 $T=224800 470995 0 90 $X=221540 $Y=470315
X1621 VSS VDD GWEN CLK 23877 1053 wen_v2 $T=208415 16605 0 0 $X=208280 $Y=15275
X1622 VSS 1 VDD CLK A[5] A[4] A[3] 1045 1046 1047 1048 1049 1050 1051 1052 xpredec1 $T=219860 111460 0 0 $X=219855 $Y=111455
X1623 VDD 1005 CLK pfet_03v3_I08 $T=234280 43425 1 0 $X=233240 $Y=41905
X1624 VDD 1006 1005 pfet_03v3_I08 $T=239670 43425 1 0 $X=238630 $Y=41905
X1625 VSS 1005 CLK nfet_03v3_I15 $T=234280 46585 1 0 $X=233600 $Y=45365
X1626 VSS 1006 1005 nfet_03v3_I15 $T=239670 46585 1 0 $X=238990 $Y=45365
X1638 VDD VSS 23266 23267 23268 23269 23270 23271 23272 23273 23943 23944 23945 23946 23947 23948 23949 23950 704 705
+ 24738 24739 24740 24741 24742 24743 24744 24745 24746 24747 24748 24749 24750 24751 24752 24753 24754 24755 24756 24757
+ ICV_31 $T=307090 180630 1 180 $X=303750 $Y=180290
X1639 VDD VSS 23274 23275 23276 23277 23278 23279 23280 23281 23943 23944 23945 23946 23947 23948 23949 23950 704 705
+ 24758 24759 24760 24761 24762 24763 24764 24765 24766 24767 24768 24769 24770 24771 24772 24773 24774 24775 24776 24777
+ ICV_31 $T=307090 216630 1 180 $X=303750 $Y=216290
X1640 VDD VSS 23282 23283 23284 23285 23286 23287 23288 23289 23943 23944 23945 23946 23947 23948 23949 23950 704 705
+ 24778 24779 24780 24781 24782 24783 24784 24785 24786 24787 24788 24789 24790 24791 24792 24793 24794 24795 24796 24797
+ ICV_31 $T=307090 252630 1 180 $X=303750 $Y=252290
X1641 VDD VSS 23290 23291 23292 23293 23294 23295 23296 23297 23943 23944 23945 23946 23947 23948 23949 23950 704 705
+ 24798 24799 24800 24801 24802 24803 24804 24805 24806 24807 24808 24809 24810 24811 24812 24813 24814 24815 24816 24817
+ ICV_31 $T=307090 288630 1 180 $X=303750 $Y=288290
X1642 VDD VSS 23298 23299 23300 23301 23302 23303 23304 23305 23943 23944 23945 23946 23947 23948 23949 23950 704 705
+ 24818 24819 24820 24821 24822 24823 24824 24825 24826 24827 24828 24829 24830 24831 24832 24833 24834 24835 24836 24837
+ ICV_31 $T=307090 324630 1 180 $X=303750 $Y=324290
X1643 VDD VSS 23306 23307 23308 23309 23310 23311 23312 23313 23943 23944 23945 23946 23947 23948 23949 23950 704 705
+ 24838 24839 24840 24841 24842 24843 24844 24845 24846 24847 24848 24849 24850 24851 24852 24853 24854 24855 24856 24857
+ ICV_31 $T=307090 360630 1 180 $X=303750 $Y=360290
X1644 VDD VSS 23314 23315 23316 23317 23318 23319 23320 23321 23943 23944 23945 23946 23947 23948 23949 23950 704 705
+ 24858 24859 24860 24861 24862 24863 24864 24865 24866 24867 24868 24869 24870 24871 24872 24873 24874 24875 24876 24877
+ ICV_31 $T=307090 396630 1 180 $X=303750 $Y=396290
X1645 VDD VSS 23322 23323 23324 23325 23326 23327 23328 23329 23943 23944 23945 23946 23947 23948 23949 23950 704 705
+ 24878 24879 24880 24881 24882 24883 24884 24885 24886 24887 24888 24889 24890 24891 24892 24893 24894 24895 24896 24897
+ ICV_31 $T=307090 432630 1 180 $X=303750 $Y=432290
X1648 614 615 VSS VDD 24074 24075 24076 24077 ICV_4 $T=415090 176130 0 0 $X=414750 $Y=175790
X1649 614 615 VSS VDD 24078 24079 24080 24081 ICV_4 $T=415090 212130 0 0 $X=414750 $Y=211790
X1650 614 615 VSS VDD 24082 24083 24084 24085 ICV_4 $T=415090 248130 0 0 $X=414750 $Y=247790
X1651 614 615 VSS VDD 24086 24087 24088 24089 ICV_4 $T=415090 284130 0 0 $X=414750 $Y=283790
X1652 614 615 VSS VDD 24090 24091 24092 24093 ICV_4 $T=415090 320130 0 0 $X=414750 $Y=319790
X1653 614 615 VSS VDD 24094 24095 24096 24097 ICV_4 $T=415090 356130 0 0 $X=414750 $Y=355790
X1654 614 615 VSS VDD 24098 24099 24100 24101 ICV_4 $T=415090 392130 0 0 $X=414750 $Y=391790
X1655 614 615 VSS VDD 24102 24103 24104 24105 ICV_4 $T=415090 428130 0 0 $X=414750 $Y=427790
.ENDS
***************************************
