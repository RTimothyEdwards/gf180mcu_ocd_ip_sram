magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal1 >>
rect -113 322 113 330
rect -113 -322 -105 322
rect 105 -322 113 322
rect -113 -330 113 -322
<< via1 >>
rect -105 -322 105 322
<< metal2 >>
rect -113 322 113 330
rect -113 -322 -105 322
rect 105 -322 113 322
rect -113 -330 113 -322
<< end >>
