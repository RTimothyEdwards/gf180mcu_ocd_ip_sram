magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< nwell >>
rect -133 -66 160 700
<< polysilicon >>
rect -14 635 41 668
rect -14 -34 41 0
use pmos_5p0431059130201_3v512x8m81  pmos_5p0431059130201_3v512x8m81_0
timestamp 1764525316
transform 1 0 -14 0 1 0
box -174 -86 230 721
<< end >>
