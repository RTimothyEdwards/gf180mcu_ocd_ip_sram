magic
tech gf180mcuD
magscale 1 10
timestamp 1763483433
<< metal1 >>
rect 2654 20538 4331 20632
rect 2632 16891 4157 17027
<< metal2 >>
rect 2831 25266 3510 36851
rect 2831 9963 3531 25266
rect 2831 1811 3531 9613
<< metal3 >>
rect 2338 25911 4138 26051
rect 2338 25784 3047 25911
rect 2338 25448 4138 25784
rect 2338 23755 4138 25160
rect 2338 22413 3531 23755
rect 2338 22214 4642 22413
rect 2338 20427 4445 21814
rect 2338 18039 3531 18429
rect 2338 17729 4445 18039
rect 2338 16952 4445 17270
rect 2338 16570 3047 16952
rect 2338 14224 4445 16130
rect 2338 11642 4445 14024
rect 2338 11036 4445 11537
rect 2338 10605 3531 11036
rect 2338 10038 4445 10605
rect 2338 8736 4445 9658
rect 2338 7319 4445 8273
rect 2338 6500 4445 6930
rect 2338 5952 3047 6500
rect 2338 5649 4445 5952
rect 2338 5234 4445 5553
rect 2338 4773 3535 5234
rect 2338 4455 4445 4773
rect 2338 4007 4445 4253
rect 2338 3611 3037 4007
rect 2338 3364 4445 3611
rect 2338 2476 4445 3176
use M2_M14310591302080_512x8m81  M2_M14310591302080_512x8m81_0
timestamp 1763476864
transform 1 0 2648 0 1 3809
box -113 -417 113 417
use M2_M14310591302080_512x8m81  M2_M14310591302080_512x8m81_1
timestamp 1763476864
transform 1 0 2648 0 1 9199
box -113 -417 113 417
use M2_M14310591302081_512x8m81  M2_M14310591302081_512x8m81_0
timestamp 1763476864
transform 1 0 2648 0 1 16761
box -113 -330 113 330
use M2_M14310591302087_512x8m81  M2_M14310591302087_512x8m81_0
timestamp 1763476864
transform 1 0 2648 0 1 25721
box -113 -243 113 243
use M2_M14310591302092_512x8m81  M2_M14310591302092_512x8m81_0
timestamp 1763476864
transform 1 0 2648 0 1 12856
box -113 -1155 113 1155
use M2_M14310591302093_512x8m81  M2_M14310591302093_512x8m81_0
timestamp 1763476864
transform 1 0 2648 0 1 6297
box -113 -634 113 634
use M2_M14310591302093_512x8m81  M2_M14310591302093_512x8m81_1
timestamp 1763476864
transform 1 0 2648 0 1 20504
box -113 -634 113 634
use M3_M24310591302042_512x8m81  M3_M24310591302042_512x8m81_0
timestamp 1763476864
transform 1 0 3189 0 1 2823
box -330 -330 330 330
use M3_M24310591302042_512x8m81  M3_M24310591302042_512x8m81_1
timestamp 1763476864
transform 1 0 3189 0 1 18060
box -330 -330 330 330
use M3_M24310591302082_512x8m81  M3_M24310591302082_512x8m81_0
timestamp 1763476864
transform 1 0 3189 0 1 5014
box -330 -547 330 547
use M3_M24310591302083_512x8m81  M3_M24310591302083_512x8m81_0
timestamp 1763476864
transform 1 0 3189 0 1 23524
box -330 -1282 330 1632
use M3_M24310591302084_512x8m81  M3_M24310591302084_512x8m81_0
timestamp 1763476864
transform 1 0 2648 0 1 12856
box -113 -1155 113 1155
use M3_M24310591302085_512x8m81  M3_M24310591302085_512x8m81_0
timestamp 1763476864
transform 1 0 2648 0 1 16921
box -113 -330 113 330
use M3_M24310591302086_512x8m81  M3_M24310591302086_512x8m81_0
timestamp 1763476864
transform 1 0 2648 0 1 6297
box -113 -634 113 634
use M3_M24310591302086_512x8m81  M3_M24310591302086_512x8m81_1
timestamp 1763476864
transform 1 0 2648 0 1 21154
box -113 -634 113 634
use M3_M24310591302088_512x8m81  M3_M24310591302088_512x8m81_0
timestamp 1763476864
transform 1 0 3189 0 1 10795
box -330 -721 330 721
use M3_M24310591302089_512x8m81  M3_M24310591302089_512x8m81_0
timestamp 1763476864
transform 1 0 2648 0 1 3809
box -113 -417 113 417
use M3_M24310591302089_512x8m81  M3_M24310591302089_512x8m81_1
timestamp 1763476864
transform 1 0 2648 0 1 9199
box -113 -417 113 417
use M3_M24310591302090_512x8m81  M3_M24310591302090_512x8m81_0
timestamp 1763476864
transform 1 0 2648 0 1 25721
box -113 -243 113 243
use M3_M24310591302091_512x8m81  M3_M24310591302091_512x8m81_0
timestamp 1763476864
transform 1 0 3189 0 1 7800
box -330 -460 330 460
use M3_M24310591302094_512x8m81  M3_M24310591302094_512x8m81_0
timestamp 1763476864
transform 1 0 3189 0 1 15177
box -330 -938 330 938
<< end >>
