magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< error_s >>
rect -173 0 -127 84
rect -13 0 33 84
rect 147 0 193 84
rect 308 0 354 84
rect 468 0 514 84
<< nwell >>
rect -133 -62 203 150
rect 204 -46 546 150
rect 204 -62 490 -46
rect -133 -66 490 -62
use pmos_5p04310591302021_3v1024x8m81  pmos_5p04310591302021_3v1024x8m81_0
timestamp 1764525316
transform 1 0 -14 0 1 0
box -258 -86 627 170
<< end >>
