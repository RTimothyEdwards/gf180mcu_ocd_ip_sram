magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -119 248 119 275
rect -119 -248 -93 248
rect 93 -248 119 248
rect -119 -275 119 -248
<< via2 >>
rect -93 -248 93 248
<< metal3 >>
rect -119 248 119 275
rect -119 -248 -93 248
rect 93 -248 119 248
rect -119 -275 119 -248
<< end >>
