magic
tech gf180mcuD
magscale 1 10
timestamp 1765833244
<< nwell >>
rect -310 -62 27 447
rect 28 -62 333 447
rect -310 -66 333 -62
rect 334 -54 653 447
rect 654 -54 983 447
rect 334 -66 983 -54
rect 984 -49 1325 447
rect 984 -65 1213 -49
rect 984 -66 1185 -65
<< polysilicon >>
rect -266 381 -211 415
rect -106 381 -50 415
rect 55 381 111 415
rect 215 381 271 415
rect 376 381 432 415
rect 536 381 592 415
rect 697 381 753 415
rect 857 381 913 415
rect 1018 381 1074 415
rect 1178 381 1234 415
rect -266 -34 -211 0
rect -106 -34 -50 0
rect 55 -34 111 0
rect 215 -34 271 0
rect 376 -34 432 0
rect 536 -34 592 0
rect 697 -34 753 0
rect 857 -34 913 0
rect 1018 -34 1074 0
rect 1178 -34 1234 0
use pmos_5p04310591302022_3v256x8m81  pmos_5p04310591302022_3v256x8m81_0
timestamp 1765833244
transform 1 0 -14 0 1 0
box -426 -86 1422 467
<< end >>
