magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< nwell >>
rect -174 -86 230 330
<< pmos >>
rect 0 0 56 244
<< pdiff >>
rect -88 231 0 244
rect -88 13 -75 231
rect -29 13 0 231
rect -88 0 0 13
rect 56 231 144 244
rect 56 13 85 231
rect 131 13 144 231
rect 56 0 144 13
<< pdiffc >>
rect -75 13 -29 231
rect 85 13 131 231
<< polysilicon >>
rect 0 244 56 288
rect 0 -44 56 0
<< metal1 >>
rect -75 231 -29 244
rect -75 0 -29 13
rect 85 231 131 244
rect 85 0 131 13
<< labels >>
flabel pdiffc -40 122 -40 122 0 FreeSans 186 0 0 0 S
flabel pdiffc 96 122 96 122 0 FreeSans 186 0 0 0 D
<< end >>
