magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nmos >>
rect 0 0 56 178
<< ndiff >>
rect -88 165 0 178
rect -88 13 -75 165
rect -29 13 0 165
rect -88 0 0 13
rect 56 165 144 178
rect 56 13 85 165
rect 131 13 144 165
rect 56 0 144 13
<< ndiffc >>
rect -75 13 -29 165
rect 85 13 131 165
<< polysilicon >>
rect 0 178 56 222
rect 0 -44 56 0
<< metal1 >>
rect -75 165 -29 178
rect -75 0 -29 13
rect 85 165 131 178
rect 85 0 131 13
<< labels >>
flabel ndiffc -40 89 -40 89 0 FreeSans 93 0 0 0 S
flabel ndiffc 96 89 96 89 0 FreeSans 93 0 0 0 D
<< end >>
