magic
tech gf180mcuD
magscale 1 10
timestamp 1763482574
<< metal2 >>
rect -75 1666 45 7039
rect 150 1428 270 6816
rect 360 1190 480 6587
rect 570 952 690 6364
rect 783 714 903 5780
rect 994 476 1114 5556
rect 1198 238 1318 5319
rect 1425 0 1545 5073
<< metal3 >>
rect -73 6920 2478 7071
rect 150 6675 2478 6826
rect 357 6430 2478 6581
rect 559 6185 2478 6335
rect 776 5661 2478 5811
rect 978 5418 2478 5569
rect 1174 5168 2478 5319
rect 1413 4924 2478 5075
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_0
timestamp 1763476864
transform -1 0 -7 0 1 1743
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_1
timestamp 1763476864
transform -1 0 219 0 1 1501
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_2
timestamp 1763476864
transform -1 0 429 0 1 1277
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_3
timestamp 1763476864
transform -1 0 640 0 1 1037
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_4
timestamp 1763476864
transform -1 0 853 0 1 803
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_5
timestamp 1763476864
transform -1 0 1064 0 1 542
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_6
timestamp 1763476864
transform -1 0 1268 0 1 317
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_7
timestamp 1763476864
transform -1 0 1485 0 1 80
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_8
timestamp 1763476864
transform -1 0 1268 0 1 5245
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_9
timestamp 1763476864
transform -1 0 1064 0 1 5495
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_10
timestamp 1763476864
transform -1 0 853 0 1 5737
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_11
timestamp 1763476864
transform -1 0 640 0 1 6261
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_12
timestamp 1763476864
transform -1 0 429 0 1 6506
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_13
timestamp 1763476864
transform -1 0 219 0 1 6747
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_14
timestamp 1763476864
transform -1 0 -7 0 1 6992
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_15
timestamp 1763476864
transform -1 0 1492 0 1 4999
box -63 -63 63 63
<< end >>
