magic
tech gf180mcuD
magscale 1 10
timestamp 1765483240
<< metal2 >>
rect 8045 119 8135 213
rect 8309 119 8400 213
rect 8573 119 8664 213
rect 8838 119 8928 213
rect 9102 119 9193 213
rect 10609 119 10699 213
rect 10873 119 10964 213
rect 11137 119 11228 213
rect 11402 119 11492 213
rect 11666 119 11757 213
rect 11930 119 12021 213
rect 12195 119 12285 213
rect 12460 119 12550 213
rect 4784 -14 4875 78
<< metal3 >>
rect 239 19374 330 19467
rect 535 19065 626 19158
rect 16350 19065 16440 19158
rect 239 18744 330 18837
rect 535 18441 626 18534
rect 16350 18441 16440 18534
rect 535 17845 626 17938
rect 16350 17845 16440 17938
rect 535 17231 626 17324
rect 16350 17231 16440 17324
rect 535 16635 626 16728
rect 16350 16635 16440 16728
rect 535 16021 626 16114
rect 16350 16011 16440 16104
rect 535 15425 626 15518
rect 16350 15425 16440 15518
rect 535 14811 626 14904
rect 16350 14801 16440 14894
rect 535 14215 626 14308
rect 16350 14215 16440 14308
rect 535 13591 626 13684
rect 16350 13591 16440 13684
rect 535 13005 626 13098
rect 16350 12995 16440 13088
rect 535 12381 626 12474
rect 16350 12381 16440 12474
rect 535 11795 626 11888
rect 16350 11785 16440 11878
rect 535 11171 626 11264
rect 16350 11171 16440 11264
rect 535 10575 626 10668
rect 16350 10575 16440 10668
rect 535 9961 626 10054
rect 16350 9951 16440 10044
rect 535 9365 626 9458
rect 16350 9365 16440 9458
rect 535 8741 626 8834
rect 16350 8741 16440 8834
rect 535 8155 626 8248
rect 16350 8155 16440 8248
rect 535 7531 626 7624
rect 16350 7531 16440 7624
rect 535 6945 626 7038
rect 16350 6935 16440 7028
rect 535 6321 626 6414
rect 16350 6311 16440 6404
rect 535 5725 626 5818
rect 16350 5725 16440 5818
rect 535 5111 626 5204
rect 16350 5101 16440 5194
rect 535 4515 626 4608
rect 16350 4515 16440 4608
rect 535 3891 626 3984
rect 16350 3891 16440 3984
rect 535 3295 626 3388
rect 16350 3305 16440 3398
rect 535 2681 626 2774
rect 16350 2681 16440 2774
rect 535 2085 626 2178
rect 16350 2095 16440 2188
rect 535 1471 626 1564
rect 16350 1471 16440 1564
rect 535 885 626 978
rect 16350 875 16440 968
rect 535 261 626 354
rect 16364 256 16456 350
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_0
timestamp 1764525316
transform 1 0 7561 0 1 166
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_1
timestamp 1764525316
transform 1 0 7561 0 1 1068
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_2
timestamp 1764525316
transform 1 0 7561 0 1 1381
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_3
timestamp 1764525316
transform 1 0 8354 0 1 15454
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_4
timestamp 1764525316
transform 1 0 8354 0 1 16085
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_5
timestamp 1764525316
transform 1 0 8354 0 1 16666
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_6
timestamp 1764525316
transform 1 0 8354 0 1 17295
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_7
timestamp 1764525316
transform 1 0 8354 0 1 17876
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_8
timestamp 1764525316
transform 1 0 8619 0 1 14241
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_9
timestamp 1764525316
transform 1 0 8354 0 1 19088
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_10
timestamp 1764525316
transform 1 0 8354 0 1 18510
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_11
timestamp 1764525316
transform 1 0 8883 0 1 5177
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_12
timestamp 1764525316
transform 1 0 8883 0 1 5754
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_13
timestamp 1764525316
transform 1 0 8883 0 1 6388
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_14
timestamp 1764525316
transform 1 0 8883 0 1 6971
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_15
timestamp 1764525316
transform 1 0 8883 0 1 7598
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_16
timestamp 1764525316
transform 1 0 8883 0 1 8181
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_17
timestamp 1764525316
transform 1 0 7561 0 1 19248
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_18
timestamp 1764525316
transform 1 0 7561 0 1 18038
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_19
timestamp 1764525316
transform 1 0 7561 0 1 16823
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_20
timestamp 1764525316
transform 1 0 7561 0 1 15610
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_21
timestamp 1764525316
transform 1 0 7561 0 1 14400
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_22
timestamp 1764525316
transform 1 0 7561 0 1 13191
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_23
timestamp 1764525316
transform 1 0 7561 0 1 11973
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_24
timestamp 1764525316
transform 1 0 7561 0 1 10763
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_25
timestamp 1764525316
transform 1 0 7561 0 1 9553
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_26
timestamp 1764525316
transform 1 0 7561 0 1 8343
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_27
timestamp 1764525316
transform 1 0 7561 0 1 7123
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_28
timestamp 1764525316
transform 1 0 7561 0 1 5913
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_29
timestamp 1764525316
transform 1 0 7561 0 1 4703
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_30
timestamp 1764525316
transform 1 0 7561 0 1 3493
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_31
timestamp 1764525316
transform 1 0 7561 0 1 2281
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_32
timestamp 1764525316
transform 1 0 8619 0 1 10026
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_33
timestamp 1764525316
transform 1 0 8619 0 1 10606
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_34
timestamp 1764525316
transform 1 0 9147 0 1 4544
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_35
timestamp 1764525316
transform 1 0 8619 0 1 11238
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_36
timestamp 1764525316
transform 1 0 8883 0 1 9394
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_37
timestamp 1764525316
transform 1 0 8883 0 1 8814
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_38
timestamp 1764525316
transform 1 0 8619 0 1 11819
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_39
timestamp 1764525316
transform 1 0 8619 0 1 12448
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_40
timestamp 1764525316
transform 1 0 8619 0 1 13029
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_41
timestamp 1764525316
transform 1 0 9147 0 1 328
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_42
timestamp 1764525316
transform 1 0 9147 0 1 906
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_43
timestamp 1764525316
transform 1 0 9147 0 1 1543
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_44
timestamp 1764525316
transform 1 0 9147 0 1 2119
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_45
timestamp 1764525316
transform 1 0 9147 0 1 2754
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_46
timestamp 1764525316
transform 1 0 9147 0 1 3331
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_47
timestamp 1764525316
transform 1 0 9147 0 1 3968
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_48
timestamp 1764525316
transform 1 0 7561 0 1 18349
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_49
timestamp 1764525316
transform 1 0 7561 0 1 17138
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_50
timestamp 1764525316
transform 1 0 7561 0 1 15923
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_51
timestamp 1764525316
transform 1 0 7561 0 1 14713
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_52
timestamp 1764525316
transform 1 0 7561 0 1 13502
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_53
timestamp 1764525316
transform 1 0 7561 0 1 12286
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_54
timestamp 1764525316
transform 1 0 7561 0 1 11076
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_55
timestamp 1764525316
transform 1 0 7561 0 1 9866
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_56
timestamp 1764525316
transform 1 0 7561 0 1 8656
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_57
timestamp 1764525316
transform 1 0 7561 0 1 7436
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_58
timestamp 1764525316
transform 1 0 7561 0 1 6226
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_59
timestamp 1764525316
transform 1 0 7561 0 1 5016
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_60
timestamp 1764525316
transform 1 0 7561 0 1 3804
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_61
timestamp 1764525316
transform 1 0 7561 0 1 2592
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_62
timestamp 1764525316
transform 1 0 8619 0 1 13658
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_63
timestamp 1764525316
transform 1 0 8354 0 1 14873
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_64
timestamp 1764525316
transform 1 0 12504 0 1 404
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_65
timestamp 1764525316
transform 1 0 12240 0 1 833
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_66
timestamp 1764525316
transform 1 0 11976 0 1 1616
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_67
timestamp 1764525316
transform 1 0 11711 0 1 2045
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_68
timestamp 1764525316
transform 1 0 11447 0 1 2827
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_69
timestamp 1764525316
transform 1 0 11183 0 1 3256
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_70
timestamp 1764525316
transform 1 0 10918 0 1 4042
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_71
timestamp 1764525316
transform 1 0 10654 0 1 4468
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_72
timestamp 1764525316
transform 1 0 10654 0 1 9315
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_73
timestamp 1764525316
transform 1 0 10654 0 1 14165
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_74
timestamp 1764525316
transform 1 0 10654 0 1 19012
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_75
timestamp 1764525316
transform 1 0 10918 0 1 8886
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_76
timestamp 1764525316
transform 1 0 10918 0 1 13736
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_77
timestamp 1764525316
transform 1 0 10918 0 1 18584
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_78
timestamp 1764525316
transform 1 0 11183 0 1 8103
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_79
timestamp 1764525316
transform 1 0 11183 0 1 12951
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_80
timestamp 1764525316
transform 1 0 11183 0 1 17803
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_81
timestamp 1764525316
transform 1 0 11447 0 1 7674
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_82
timestamp 1764525316
transform 1 0 11447 0 1 12522
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_83
timestamp 1764525316
transform 1 0 11447 0 1 17374
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_84
timestamp 1764525316
transform 1 0 11711 0 1 6891
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_85
timestamp 1764525316
transform 1 0 11711 0 1 11741
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_86
timestamp 1764525316
transform 1 0 11711 0 1 16587
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_87
timestamp 1764525316
transform 1 0 11976 0 1 6463
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_88
timestamp 1764525316
transform 1 0 11976 0 1 11312
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_89
timestamp 1764525316
transform 1 0 11976 0 1 16156
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_90
timestamp 1764525316
transform 1 0 12240 0 1 5681
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_91
timestamp 1764525316
transform 1 0 12240 0 1 10529
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_92
timestamp 1764525316
transform 1 0 12240 0 1 15375
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_93
timestamp 1764525316
transform 1 0 12504 0 1 5252
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_94
timestamp 1764525316
transform 1 0 12504 0 1 10100
box -44 -46 44 46
use M2_M1$$202394668_3v1024x8m81  M2_M1$$202394668_3v1024x8m81_95
timestamp 1764525316
transform 1 0 12504 0 1 14946
box -44 -46 44 46
use xdec8_3v1024x8m81  xdec8_3v1024x8m81_0
timestamp 1764692000
transform 1 0 0 0 1 14544
box 230 -159 16952 5031
use xdec8_3v1024x8m81  xdec8_3v1024x8m81_1
timestamp 1764692000
transform 1 0 0 0 1 0
box 230 -159 16952 5031
use xdec8_3v1024x8m81  xdec8_3v1024x8m81_2
timestamp 1764692000
transform 1 0 0 0 1 4848
box 230 -159 16952 5031
use xdec8_3v1024x8m81  xdec8_3v1024x8m81_3
timestamp 1764692000
transform 1 0 0 0 1 9696
box 230 -159 16952 5031
<< labels >>
rlabel metal3 s 581 308 581 308 4 LWL[0]
port 12 nsew
rlabel metal3 s 16396 308 16396 308 4 RWL[0]
port 26 nsew
rlabel metal2 s 11976 166 11976 166 4 xa[2]
port 67 nsew
rlabel metal2 s 4830 31 4830 31 4 men
port 68 nsew
rlabel metal2 s 12504 166 12504 166 4 xa[0]
port 69 nsew
rlabel metal2 s 11711 166 11711 166 4 xa[3]
port 70 nsew
rlabel metal2 s 11447 166 11447 166 4 xa[4]
port 71 nsew
rlabel metal2 s 11183 166 11183 166 4 xa[5]
port 72 nsew
rlabel metal2 s 10918 166 10918 166 4 xa[6]
port 73 nsew
rlabel metal2 s 10654 166 10654 166 4 xa[7]
port 74 nsew
rlabel metal2 s 8354 166 8354 166 4 xb[3]
port 75 nsew
rlabel metal2 s 8619 166 8619 166 4 xb[2]
port 76 nsew
rlabel metal2 s 8883 166 8883 166 4 xb[1]
port 77 nsew
rlabel metal2 s 9147 166 9147 166 4 xb[0]
port 78 nsew
rlabel metal2 s 8090 166 8090 166 4 xc
port 79 nsew
rlabel metal2 s 12240 166 12240 166 4 xa[1]
port 80 nsew
rlabel metal3 s 16396 922 16396 922 4 RWL[1]
port 25 nsew
rlabel metal3 s 16396 1518 16396 1518 4 RWL[2]
port 27 nsew
rlabel metal3 s 16396 2142 16396 2142 4 RWL[3]
port 24 nsew
rlabel metal3 s 16396 2728 16396 2728 4 RWL[4]
port 37 nsew
rlabel metal3 s 16396 3352 16396 3352 4 RWL[5]
port 23 nsew
rlabel metal3 s 16396 3938 16396 3938 4 RWL[6]
port 38 nsew
rlabel metal3 s 16396 4562 16396 4562 4 RWL[7]
port 22 nsew
rlabel metal3 s 16396 5148 16396 5148 4 RWL[8]
port 21 nsew
rlabel metal3 s 16396 5772 16396 5772 4 RWL[9]
port 20 nsew
rlabel metal3 s 16396 6358 16396 6358 4 RWL[10]
port 19 nsew
rlabel metal3 s 16396 6982 16396 6982 4 RWL[11]
port 18 nsew
rlabel metal3 s 16396 7578 16396 7578 4 RWL[12]
port 9 nsew
rlabel metal3 s 16396 8202 16396 8202 4 RWL[13]
port 8 nsew
rlabel metal3 s 16396 8788 16396 8788 4 RWL[14]
port 7 nsew
rlabel metal3 s 16396 9412 16396 9412 4 RWL[15]
port 6 nsew
rlabel metal3 s 16396 9998 16396 9998 4 RWL[16]
port 5 nsew
rlabel metal3 s 16396 10622 16396 10622 4 RWL[17]
port 4 nsew
rlabel metal3 s 16396 11218 16396 11218 4 RWL[18]
port 3 nsew
rlabel metal3 s 16396 11832 16396 11832 4 RWL[19]
port 66 nsew
rlabel metal3 s 16396 12428 16396 12428 4 RWL[20]
port 49 nsew
rlabel metal3 s 16396 13042 16396 13042 4 RWL[21]
port 50 nsew
rlabel metal3 s 16396 13638 16396 13638 4 RWL[22]
port 51 nsew
rlabel metal3 s 16396 14262 16396 14262 4 RWL[23]
port 52 nsew
rlabel metal3 s 16396 14848 16396 14848 4 RWL[24]
port 53 nsew
rlabel metal3 s 16396 15472 16396 15472 4 RWL[25]
port 54 nsew
rlabel metal3 s 16396 16058 16396 16058 4 RWL[26]
port 55 nsew
rlabel metal3 s 16396 16682 16396 16682 4 RWL[27]
port 56 nsew
rlabel metal3 s 16396 17278 16396 17278 4 RWL[28]
port 57 nsew
rlabel metal3 s 16396 17892 16396 17892 4 RWL[29]
port 58 nsew
rlabel metal3 s 16396 18488 16396 18488 4 RWL[30]
port 59 nsew
rlabel metal3 s 16396 19112 16396 19112 4 RWL[31]
port 60 nsew
rlabel metal3 s 581 932 581 932 4 LWL[1]
port 13 nsew
rlabel metal3 s 581 1518 581 1518 4 LWL[2]
port 14 nsew
rlabel metal3 s 581 2132 581 2132 4 LWL[3]
port 15 nsew
rlabel metal3 s 581 2728 581 2728 4 LWL[4]
port 16 nsew
rlabel metal3 s 581 3342 581 3342 4 LWL[5]
port 17 nsew
rlabel metal3 s 581 3938 581 3938 4 LWL[6]
port 1 nsew
rlabel metal3 s 581 4562 581 4562 4 LWL[7]
port 2 nsew
rlabel metal3 s 581 5158 581 5158 4 LWL[8]
port 11 nsew
rlabel metal3 s 581 5772 581 5772 4 LWL[9]
port 10 nsew
rlabel metal3 s 581 6368 581 6368 4 LWL[10]
port 36 nsew
rlabel metal3 s 581 6992 581 6992 4 LWL[11]
port 35 nsew
rlabel metal3 s 581 7578 581 7578 4 LWL[12]
port 34 nsew
rlabel metal3 s 581 8202 581 8202 4 LWL[13]
port 33 nsew
rlabel metal3 s 581 8788 581 8788 4 LWL[14]
port 32 nsew
rlabel metal3 s 581 9412 581 9412 4 LWL[15]
port 31 nsew
rlabel metal3 s 581 10008 581 10008 4 LWL[16]
port 30 nsew
rlabel metal3 s 581 10622 581 10622 4 LWL[17]
port 29 nsew
rlabel metal3 s 581 11218 581 11218 4 LWL[18]
port 28 nsew
rlabel metal3 s 581 11842 581 11842 4 LWL[19]
port 48 nsew
rlabel metal3 s 581 12428 581 12428 4 LWL[20]
port 47 nsew
rlabel metal3 s 581 13052 581 13052 4 LWL[21]
port 46 nsew
rlabel metal3 s 581 13638 581 13638 4 LWL[22]
port 45 nsew
rlabel metal3 s 581 14262 581 14262 4 LWL[23]
port 44 nsew
rlabel metal3 s 581 14858 581 14858 4 LWL[24]
port 43 nsew
rlabel metal3 s 581 15472 581 15472 4 LWL[25]
port 42 nsew
rlabel metal3 s 581 16068 581 16068 4 LWL[26]
port 41 nsew
rlabel metal3 s 581 16682 581 16682 4 LWL[27]
port 40 nsew
rlabel metal3 s 581 17278 581 17278 4 LWL[28]
port 39 nsew
rlabel metal3 s 581 17892 581 17892 4 LWL[29]
port 63 nsew
rlabel metal3 s 581 18488 581 18488 4 LWL[30]
port 62 nsew
rlabel metal3 s 581 19112 581 19112 4 LWL[31]
port 61 nsew
rlabel metal3 s 284 19421 284 19421 4 vdd
port 64 nsew
rlabel metal3 s 284 18791 284 18791 4 vss
port 65 nsew
<< end >>
