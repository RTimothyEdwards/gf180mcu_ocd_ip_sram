magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< error_p >>
rect -75 0 -29 84
rect 141 0 187 84
<< nwell >>
rect -174 -86 286 170
<< pmos >>
rect 0 0 112 84
<< pdiff >>
rect -88 71 0 84
rect -88 13 -75 71
rect -29 13 0 71
rect -88 0 0 13
rect 112 71 200 84
rect 112 13 141 71
rect 187 13 200 71
rect 112 0 200 13
<< pdiffc >>
rect -75 13 -29 71
rect 141 13 187 71
<< polysilicon >>
rect 0 84 112 128
rect 0 -44 112 0
<< metal1 >>
rect -75 71 -29 84
rect -75 0 -29 13
rect 141 71 187 84
rect 141 0 187 13
<< labels >>
flabel pdiffc -40 42 -40 42 0 FreeSans 186 0 0 0 S
flabel pdiffc 152 42 152 42 0 FreeSans 186 0 0 0 D
<< end >>
