magic
tech gf180mcuD
magscale 1 10
timestamp 1764626446
<< nwell >>
rect 30 512 570 797
<< pwell >>
rect 82 89 518 512
<< sramnfet >>
rect 192 342 248 432
rect 352 342 408 432
rect 110 178 166 250
rect 434 178 490 250
<< srampfet >>
rect 192 592 248 648
rect 352 592 408 648
<< sramndiff >>
rect 110 424 192 432
rect 110 378 117 424
rect 163 378 192 424
rect 110 342 192 378
rect 248 342 352 432
rect 408 424 490 432
rect 408 378 437 424
rect 483 378 490 424
rect 408 342 490 378
rect 110 250 166 342
rect 270 327 330 342
rect 270 281 277 327
rect 323 281 330 327
rect 270 270 330 281
rect 434 250 490 342
rect 110 156 166 178
rect 434 156 490 178
rect 110 149 170 156
rect 110 103 117 149
rect 163 103 170 149
rect 110 96 170 103
rect 430 149 490 156
rect 430 103 437 149
rect 483 103 490 149
rect 430 96 490 103
<< srampdiff >>
rect 270 755 330 766
rect 270 709 277 755
rect 323 709 330 755
rect 110 648 170 654
rect 270 648 330 709
rect 430 648 490 654
rect 110 647 192 648
rect 110 601 117 647
rect 163 601 192 647
rect 110 592 192 601
rect 248 592 352 648
rect 408 647 490 648
rect 408 601 437 647
rect 483 601 490 647
rect 408 592 490 601
<< sramndc >>
rect 117 378 163 424
rect 437 378 483 424
rect 277 281 323 327
rect 117 103 163 149
rect 437 103 483 149
<< srampdc >>
rect 277 709 323 755
rect 117 601 163 647
rect 437 601 483 647
<< polysilicon >>
rect 192 648 248 692
rect 352 648 408 692
rect 192 524 248 592
rect 352 572 408 592
rect 329 559 408 572
rect 192 511 271 524
rect 192 465 212 511
rect 258 465 271 511
rect 329 513 342 559
rect 388 513 408 559
rect 329 500 408 513
rect 192 452 271 465
rect 192 432 248 452
rect 352 432 408 500
rect 192 298 248 342
rect 352 298 408 342
rect 62 178 110 250
rect 166 178 434 250
rect 490 178 538 250
<< polycontact >>
rect 212 465 258 511
rect 342 513 388 559
<< metal1 >>
rect 82 755 518 760
rect 82 709 277 755
rect 323 709 518 755
rect 82 704 518 709
rect 114 647 163 657
rect 434 647 486 658
rect 114 601 117 647
rect 163 601 388 647
rect 434 601 437 647
rect 483 601 486 647
rect 114 597 388 601
rect 114 424 166 597
rect 331 559 388 597
rect 114 378 117 424
rect 163 378 166 424
rect 212 511 268 530
rect 258 465 268 511
rect 331 513 342 559
rect 331 494 388 513
rect 212 448 268 465
rect 435 448 486 601
rect 212 424 486 448
rect 212 402 437 424
rect 114 367 166 378
rect 434 378 437 402
rect 483 378 486 424
rect 434 367 486 378
rect 252 327 348 356
rect 252 321 277 327
rect 82 281 277 321
rect 323 321 348 327
rect 323 281 518 321
rect 82 199 518 281
rect 106 149 164 152
rect 106 103 117 149
rect 163 103 164 149
rect 106 100 164 103
rect 216 100 258 152
rect 342 100 384 152
rect 436 149 494 152
rect 436 103 437 149
rect 483 103 494 149
rect 436 100 494 103
<< via1 >>
rect 164 100 216 152
rect 384 100 436 152
<< metal2 >>
rect 134 152 254 771
rect 134 100 164 152
rect 216 100 254 152
rect 134 89 254 100
rect 346 152 466 771
rect 346 100 384 152
rect 436 100 466 152
rect 346 89 466 100
<< metal3 >>
rect 82 330 518 690
<< properties >>
string FIXED_BBOX 82 126 518 732
string MASKHINTS_SRAMDEF 24 89 576 797
<< end >>
