magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal1 >>
rect -119 247 119 275
rect -119 -247 -92 247
rect 92 -247 119 247
rect -119 -275 119 -247
<< via1 >>
rect -92 -247 92 247
<< metal2 >>
rect -118 247 119 275
rect -118 -247 -92 247
rect 92 -247 119 247
rect -118 -275 119 -247
<< end >>
