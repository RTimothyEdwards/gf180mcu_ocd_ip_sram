magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< nwell >>
rect -174 -86 230 1610
<< pmos >>
rect 0 0 56 1524
<< pdiff >>
rect -88 1511 0 1524
rect -88 13 -75 1511
rect -29 13 0 1511
rect -88 0 0 13
rect 56 1511 144 1524
rect 56 13 85 1511
rect 131 13 144 1511
rect 56 0 144 13
<< pdiffc >>
rect -75 13 -29 1511
rect 85 13 131 1511
<< polysilicon >>
rect 0 1524 56 1568
rect 0 -44 56 0
<< metal1 >>
rect -75 1511 -29 1524
rect -75 0 -29 13
rect 85 1511 131 1524
rect 85 0 131 13
<< labels >>
flabel pdiffc -40 762 -40 762 0 FreeSans 186 0 0 0 S
flabel pdiffc 96 762 96 762 0 FreeSans 186 0 0 0 D
<< end >>
