magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< psubdiff >>
rect -54 23 54 56
rect -54 -23 -23 23
rect 23 -23 54 23
rect -54 -56 54 -23
<< psubdiffcont >>
rect -23 -23 23 23
<< metal1 >>
rect -40 23 40 42
rect -40 -23 -23 23
rect 23 -23 40 23
rect -40 -42 40 -23
<< end >>
