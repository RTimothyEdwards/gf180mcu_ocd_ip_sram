magic
tech gf180mcuD
magscale 1 10
timestamp 1764700137
<< error_p >>
rect -35 28 35 35
rect -35 -28 -28 28
rect -35 -35 35 -28
<< metal2 >>
rect -35 28 35 35
rect -35 -28 -28 28
rect 28 -28 35 28
rect -35 -35 35 -28
<< via2 >>
rect -28 -28 28 28
<< metal3 >>
rect -35 28 35 35
rect -35 -28 -28 28
rect 28 -28 35 28
rect -35 -35 35 -28
<< end >>
