magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect 300 724 389 948
rect 300 115 389 129
<< polysilicon >>
rect 525 4851 580 4964
rect 525 4840 589 4851
rect 533 3975 589 4840
rect 895 4169 949 5016
<< metal1 >>
rect 226 4991 529 5901
rect 605 4929 686 5034
rect 605 4845 901 4929
rect 193 2291 529 4755
rect 605 3850 686 4845
rect 978 3839 1024 5115
rect -74 2154 1232 2219
rect -74 2013 1232 2078
rect -74 1871 1232 1936
rect -74 1730 1232 1795
<< metal2 >>
rect 294 5288 529 5838
rect 294 951 385 4934
rect 800 989 890 2374
rect 1143 1130 1233 2557
rect 800 896 1233 989
<< metal3 >>
rect 0 5263 1276 5898
rect -4 3120 1179 5026
rect 4 2538 1233 2632
rect 10 2281 1270 2374
use alatch_512x8m81  alatch_512x8m81_0
timestamp 1763476864
transform 1 0 49 0 1 -442
box -63 0 1196 2077
use M1_NWELL11_512x8m81  M1_NWELL11_512x8m81_0
timestamp 1763476864
transform 1 0 233 0 1 3489
box -154 -1302 154 1302
use M1_POLY2$$46559276_512x8m81  M1_POLY2$$46559276_512x8m81_0
timestamp 1763476864
transform 1 0 805 0 1 4887
box -123 -48 123 48
use M1_POLY2$$46559276_512x8m81  M1_POLY2$$46559276_512x8m81_1
timestamp 1763476864
transform 1 0 448 0 1 4887
box -123 -48 123 48
use M1_PSUB$$47335468_512x8m81  M1_PSUB$$47335468_512x8m81_0
timestamp 1763476864
transform 1 0 276 0 1 5473
box -55 -400 56 400
use M2_M1$$34864172_512x8m81  M2_M1$$34864172_512x8m81_0
timestamp 1763476864
transform 1 0 413 0 1 4887
box -119 -46 119 46
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1763476864
transform 1 0 339 0 1 1042
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_1
timestamp 1763476864
transform 1 0 645 0 1 2413
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_2
timestamp 1763476864
transform 1 0 1005 0 1 3048
box -43 -122 43 122
use M2_M1$$43376684_512x8m81  M2_M1$$43376684_512x8m81_0
timestamp 1763476864
transform 1 0 853 0 1 4067
box -44 -579 44 579
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_0
timestamp 1763476864
transform 1 0 339 0 1 5563
box -44 -275 44 275
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_1
timestamp 1763476864
transform 1 0 484 0 1 5563
box -44 -275 44 275
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_2
timestamp 1763476864
transform 1 0 848 0 1 5547
box -44 -275 44 275
use M2_M1$$47500332_512x8m81  M2_M1$$47500332_512x8m81_0
timestamp 1763476864
transform 1 0 493 0 1 3908
box -44 -732 44 732
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_0
timestamp 1763476864
transform 1 0 1188 0 1 2585
box -44 -123 44 123
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_1
timestamp 1763476864
transform 1 0 845 0 1 2251
box -44 -123 44 123
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_0
timestamp 1763476864
transform 1 0 339 0 1 5563
box -45 -275 45 275
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_1
timestamp 1763476864
transform 1 0 484 0 1 5563
box -45 -275 45 275
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_2
timestamp 1763476864
transform 1 0 848 0 1 5547
box -45 -275 45 275
use M3_M2$$47644716_512x8m81  M3_M2$$47644716_512x8m81_0
timestamp 1763476864
transform 1 0 493 0 1 3908
box -45 -732 45 732
use M3_M2$$47645740_512x8m81  M3_M2$$47645740_512x8m81_0
timestamp 1763476864
transform 1 0 853 0 1 4067
box -45 -579 45 579
use nmos_1p2$$47502380_512x8m81  nmos_1p2$$47502380_512x8m81_0
timestamp 1763476864
transform 1 0 907 0 1 5041
box -102 -44 130 531
use nmos_5p04310591302066_512x8m81  nmos_5p04310591302066_512x8m81_0
timestamp 1763476864
transform 1 0 525 0 1 4986
box -88 -44 144 701
use pmos_1p2$$47503404_512x8m81  pmos_1p2$$47503404_512x8m81_0
timestamp 1763476864
transform 1 0 547 0 1 2284
box -188 -86 216 1737
use pmos_1p2$$47504428_512x8m81  pmos_1p2$$47504428_512x8m81_0
timestamp 1763476864
transform 1 0 907 0 1 2919
box -188 -86 216 1314
<< end >>
