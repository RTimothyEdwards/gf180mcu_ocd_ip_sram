magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< nwell >>
rect -426 -86 1422 467
<< pmos >>
rect -252 0 -196 381
rect -92 0 -36 381
rect 69 0 125 381
rect 229 0 285 381
rect 390 0 446 381
rect 550 0 606 381
rect 711 0 767 381
rect 871 0 927 381
rect 1032 0 1088 381
rect 1192 0 1248 381
<< pdiff >>
rect -340 368 -252 381
rect -340 13 -327 368
rect -281 13 -252 368
rect -340 0 -252 13
rect -196 368 -92 381
rect -196 13 -167 368
rect -121 13 -92 368
rect -196 0 -92 13
rect -36 368 69 381
rect -36 13 -7 368
rect 39 13 69 368
rect -36 0 69 13
rect 125 368 229 381
rect 125 13 154 368
rect 200 13 229 368
rect 125 0 229 13
rect 285 368 390 381
rect 285 13 314 368
rect 360 13 390 368
rect 285 0 390 13
rect 446 368 550 381
rect 446 13 475 368
rect 521 13 550 368
rect 446 0 550 13
rect 606 368 711 381
rect 606 13 635 368
rect 681 13 711 368
rect 606 0 711 13
rect 767 368 871 381
rect 767 13 796 368
rect 842 13 871 368
rect 767 0 871 13
rect 927 368 1032 381
rect 927 13 956 368
rect 1002 13 1032 368
rect 927 0 1032 13
rect 1088 368 1192 381
rect 1088 13 1117 368
rect 1163 13 1192 368
rect 1088 0 1192 13
rect 1248 368 1336 381
rect 1248 13 1277 368
rect 1323 13 1336 368
rect 1248 0 1336 13
<< pdiffc >>
rect -327 13 -281 368
rect -167 13 -121 368
rect -7 13 39 368
rect 154 13 200 368
rect 314 13 360 368
rect 475 13 521 368
rect 635 13 681 368
rect 796 13 842 368
rect 956 13 1002 368
rect 1117 13 1163 368
rect 1277 13 1323 368
<< polysilicon >>
rect -252 381 -196 426
rect -92 381 -36 426
rect 69 381 125 426
rect 229 381 285 426
rect 390 381 446 426
rect 550 381 606 426
rect 711 381 767 426
rect 871 381 927 426
rect 1032 381 1088 426
rect 1192 381 1248 426
rect -252 -44 -196 0
rect -92 -44 -36 0
rect 69 -44 125 0
rect 229 -44 285 0
rect 390 -44 446 0
rect 550 -44 606 0
rect 711 -44 767 0
rect 871 -44 927 0
rect 1032 -44 1088 0
rect 1192 -44 1248 0
<< metal1 >>
rect -327 368 -281 381
rect -327 0 -281 13
rect -167 368 -121 381
rect -167 0 -121 13
rect -7 368 39 381
rect -7 0 39 13
rect 154 368 200 381
rect 154 0 200 13
rect 314 368 360 381
rect 314 0 360 13
rect 475 368 521 381
rect 475 0 521 13
rect 635 368 681 381
rect 635 0 681 13
rect 796 368 842 381
rect 796 0 842 13
rect 956 368 1002 381
rect 956 0 1002 13
rect 1117 368 1163 381
rect 1117 0 1163 13
rect 1277 368 1323 381
rect 1277 0 1323 13
<< labels >>
flabel pdiffc 498 190 498 190 0 FreeSans 186 0 0 0 D
flabel pdiffc 349 190 349 190 0 FreeSans 186 0 0 0 S
flabel pdiffc 189 190 189 190 0 FreeSans 186 0 0 0 D
flabel pdiffc 28 190 28 190 0 FreeSans 186 0 0 0 S
flabel pdiffc -132 190 -132 190 0 FreeSans 186 0 0 0 D
flabel pdiffc -292 190 -292 190 0 FreeSans 186 0 0 0 S
flabel pdiffc 807 190 807 190 0 FreeSans 186 0 0 0 D
flabel pdiffc 1128 190 1128 190 0 FreeSans 186 0 0 0 D
flabel pdiffc 645 190 645 190 0 FreeSans 186 0 0 0 S
flabel pdiffc 967 190 967 190 0 FreeSans 186 0 0 0 S
flabel pdiffc 1288 190 1288 190 0 FreeSans 186 0 0 0 S
<< end >>
