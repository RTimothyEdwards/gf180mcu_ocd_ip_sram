magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal1 >>
rect -1299 94 1299 123
rect -1299 -94 -1272 94
rect 1272 -94 1299 94
rect -1299 -123 1299 -94
<< via1 >>
rect -1272 -94 1272 94
<< metal2 >>
rect -1299 94 1299 122
rect -1299 -94 -1272 94
rect 1272 -94 1299 94
rect -1299 -123 1299 -94
<< end >>
