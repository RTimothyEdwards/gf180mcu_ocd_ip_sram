magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< error_p >>
rect -284 -54 284 53
<< nsubdiff >>
rect -284 23 284 53
rect -284 -23 -252 23
rect 252 -23 284 23
rect -284 -54 284 -23
<< nsubdiffcont >>
rect -252 -23 252 23
<< metal1 >>
rect -270 23 270 40
rect -270 -23 -252 23
rect 252 -23 270 23
rect -270 -40 270 -23
<< end >>
