magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -118 181 119 198
rect -118 -181 -102 181
rect 102 -181 119 181
rect -118 -198 119 -181
<< via2 >>
rect -102 -181 102 181
<< metal3 >>
rect -119 181 119 198
rect -119 -181 -102 181
rect 102 -181 119 181
rect -119 -198 119 -181
<< end >>
