magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< polysilicon >>
rect -67 23 67 47
rect -67 -23 -23 23
rect 23 -23 67 23
rect -67 -48 67 -23
<< polycontact >>
rect -23 -23 23 23
<< metal1 >>
rect -40 23 39 41
rect -40 -23 -23 23
rect 23 -23 39 23
rect -40 -42 39 -23
<< end >>
