magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -35 497 35 504
rect -35 -497 -28 497
rect 28 -497 35 497
rect -35 -504 35 -497
<< via2 >>
rect -28 -497 28 497
<< metal3 >>
rect -35 497 35 504
rect -35 -497 -28 497
rect 28 -497 35 497
rect -35 -504 35 -497
<< end >>
