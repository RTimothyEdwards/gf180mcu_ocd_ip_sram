magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal1 >>
rect 9103 4662 9184 4746
rect 9103 4499 9184 4583
rect 10517 4449 10567 4501
rect 9103 3926 9184 4010
rect 10517 4008 10567 4060
rect 9103 3764 9184 3848
rect 9103 3452 9184 3536
rect 9103 3289 9184 3373
rect 10517 3239 10567 3291
rect 10517 2798 10567 2850
rect 9103 2706 9184 2790
rect 9103 2544 9184 2628
rect 9103 2242 9184 2326
rect 9103 2079 9184 2163
rect 10517 2029 10567 2081
rect 9103 1496 9184 1580
rect 10517 1578 10567 1630
rect 9103 1334 9184 1418
rect 9103 1022 9184 1106
rect 9103 859 9184 943
rect 10517 809 10567 861
rect 10517 378 10567 430
rect 9103 286 9184 370
rect 9103 124 9184 208
<< metal2 >>
rect 4785 -14 4876 78
<< metal3 >>
rect 244 4820 334 4913
rect 550 4535 613 4600
rect 16365 4525 16427 4590
rect 244 4190 334 4283
rect 550 3919 613 3984
rect 16365 3909 16427 3974
rect 550 3313 613 3378
rect 16365 3313 16427 3378
rect 550 2699 613 2764
rect 16365 2699 16427 2764
rect 550 2103 613 2168
rect 16365 2113 16427 2178
rect 550 1489 613 1554
rect 16365 1489 16427 1554
rect 550 888 613 953
rect 16365 898 16427 963
rect 550 289 613 354
use xdec_3v256x8m81  xdec_3v256x8m81_0
timestamp 1763766357
transform 1 0 0 0 -1 4266
box 230 -156 16952 789
use xdec_3v256x8m81  xdec_3v256x8m81_1
timestamp 1763766357
transform 1 0 0 0 -1 3054
box 230 -156 16952 789
use xdec_3v256x8m81  xdec_3v256x8m81_2
timestamp 1763766357
transform 1 0 0 0 -1 1842
box 230 -156 16952 789
use xdec_3v256x8m81  xdec_3v256x8m81_3
timestamp 1763766357
transform 1 0 0 0 -1 630
box 230 -156 16952 789
use xdec_3v256x8m81  xdec_3v256x8m81_4
timestamp 1763766357
transform 1 0 0 0 1 4242
box 230 -156 16952 789
use xdec_3v256x8m81  xdec_3v256x8m81_5
timestamp 1763766357
transform 1 0 0 0 1 3030
box 230 -156 16952 789
use xdec_3v256x8m81  xdec_3v256x8m81_6
timestamp 1763766357
transform 1 0 0 0 1 1818
box 230 -156 16952 789
use xdec_3v256x8m81  xdec_3v256x8m81_7
timestamp 1763766357
transform 1 0 0 0 1 606
box 230 -156 16952 789
<< labels >>
rlabel metal3 s 16396 322 16396 322 4 RWL[0]
port 1 nsew
rlabel metal3 s 581 322 581 322 4 LWL[0]
port 14 nsew
rlabel metal2 s 4830 31 4830 31 4 men
port 19 nsew
rlabel metal1 s 9144 166 9144 166 4 xc
port 20 nsew
rlabel metal1 s 10542 404 10542 404 4 xa[0]
port 27 nsew
rlabel metal1 s 9144 328 9144 328 4 xb
port 21 nsew
rlabel metal3 s 289 4867 289 4867 4 vdd
port 17 nsew
rlabel metal3 s 289 4237 289 4237 4 vss
port 16 nsew
rlabel metal3 s 581 920 581 920 4 LWL[1]
port 11 nsew
rlabel metal3 s 581 1522 581 1522 4 LWL[2]
port 4 nsew
rlabel metal3 s 581 2136 581 2136 4 LWL[3]
port 15 nsew
rlabel metal3 s 581 2732 581 2732 4 LWL[4]
port 3 nsew
rlabel metal3 s 581 3346 581 3346 4 LWL[5]
port 2 nsew
rlabel metal3 s 581 3952 581 3952 4 LWL[6]
port 13 nsew
rlabel metal3 s 581 4568 581 4568 4 LWL[7]
port 12 nsew
rlabel metal3 s 16396 930 16396 930 4 RWL[1]
port 8 nsew
rlabel metal3 s 16396 1522 16396 1522 4 RWL[2]
port 7 nsew
rlabel metal3 s 16396 2146 16396 2146 4 RWL[3]
port 18 nsew
rlabel metal3 s 16396 2732 16396 2732 4 RWL[4]
port 6 nsew
rlabel metal3 s 16396 3346 16396 3346 4 RWL[5]
port 5 nsew
rlabel metal3 s 16396 3942 16396 3942 4 RWL[6]
port 10 nsew
rlabel metal3 s 16396 4558 16396 4558 4 RWL[7]
port 9 nsew
rlabel metal1 s 10542 835 10542 835 4 xa[1]
port 28 nsew
rlabel metal1 s 10542 1604 10542 1604 4 xa[2]
port 29 nsew
rlabel metal1 s 10542 2055 10542 2055 4 xa[3]
port 23 nsew
rlabel metal1 s 10542 2824 10542 2824 4 xa[4]
port 22 nsew
rlabel metal1 s 10542 3265 10542 3265 4 xa[5]
port 24 nsew
rlabel metal1 s 10542 4034 10542 4034 4 xa[6]
port 25 nsew
rlabel metal1 s 10542 4475 10542 4475 4 xa[7]
port 26 nsew
rlabel metal1 s 9144 901 9144 901 4 xb
port 21 nsew
rlabel metal1 s 9144 1064 9144 1064 4 xc
port 20 nsew
rlabel metal1 s 9144 1376 9144 1376 4 xc
port 20 nsew
rlabel metal1 s 9144 1538 9144 1538 4 xb
port 21 nsew
rlabel metal1 s 9144 2284 9144 2284 4 xc
port 20 nsew
rlabel metal1 s 9144 2121 9144 2121 4 xb
port 21 nsew
rlabel metal1 s 9144 2586 9144 2586 4 xc
port 20 nsew
rlabel metal1 s 9144 2748 9144 2748 4 xb
port 21 nsew
rlabel metal1 s 9144 3494 9144 3494 4 xc
port 20 nsew
rlabel metal1 s 9144 3331 9144 3331 4 xb
port 21 nsew
rlabel metal1 s 9144 3806 9144 3806 4 xc
port 20 nsew
rlabel metal1 s 9144 3968 9144 3968 4 xb
port 21 nsew
rlabel metal1 s 9144 4704 9144 4704 4 xc
port 20 nsew
rlabel metal1 s 9144 4541 9144 4541 4 xb
port 21 nsew
<< end >>
