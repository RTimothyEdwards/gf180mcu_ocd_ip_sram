magic
tech gf180mcuD
magscale 1 10
timestamp 1763486358
<< nwell >>
rect 225 20099 4028 20386
rect 225 18646 3458 20099
rect 225 17041 4028 18646
rect 1013 6563 1054 6600
rect 1576 6561 1612 6580
<< metal1 >>
rect 232 18911 375 18962
rect 3740 7388 3806 8070
rect 1918 6452 1976 6668
rect 2391 5599 2534 5814
rect 1269 1054 1350 1164
rect 1677 974 1736 1049
rect 1838 974 1888 1040
rect 2342 974 2389 1040
rect 1834 599 1918 731
rect 2356 599 2426 731
<< metal2 >>
rect 148 18906 264 18974
rect 26 11631 91 18824
rect 148 11519 215 18906
rect 271 11631 337 18824
rect 425 11920 488 13538
rect 1276 11987 1339 13506
rect 2199 11987 2261 13496
rect 3100 11987 3163 13490
rect 3872 11842 3935 13509
rect 3531 11774 3935 11842
rect 148 11451 439 11519
rect 660 7468 1341 7527
rect 1450 7519 1516 11520
rect 324 340 389 6238
rect 581 5777 648 6558
rect 581 5683 810 5777
rect 744 4481 810 5683
rect 1282 5728 1341 7468
rect 1579 5802 1645 11519
rect 1708 7519 1774 11520
rect 2963 6181 3028 6302
rect 3284 6269 3350 6302
rect 3284 6201 3535 6269
rect 2963 6113 3104 6181
rect 3469 6050 3535 6201
rect 1282 5669 1405 5728
rect 1579 5720 1992 5802
rect 591 4407 810 4481
rect 591 1393 658 4407
rect 1047 4356 1113 5012
rect 1346 4574 1405 5669
rect 935 4277 1113 4356
rect 1296 4514 1405 4574
rect 935 3765 1001 4277
rect 915 3691 1001 3765
rect 915 1331 981 3691
rect 1296 1644 1355 4514
rect 1608 4437 1647 4441
rect 1589 3832 1647 4437
rect 1925 3867 1992 5720
rect 3740 4570 3806 7410
rect 3059 4476 3303 4570
rect 3245 4214 3303 4476
rect 3585 4476 3806 4570
rect 3585 4214 3644 4476
rect 1495 3793 1647 3832
rect 1726 3803 1992 3867
rect 1726 3616 1803 3803
rect 1579 3555 1803 3616
rect 1579 2667 1645 3555
rect 1296 1585 1375 1644
rect 637 233 704 1296
rect 915 1258 1001 1331
rect 935 340 1001 1258
rect 1316 1034 1375 1585
rect 1316 975 1421 1034
rect 1362 278 1421 975
rect 1362 211 1741 278
rect 1682 -975 1741 211
rect 1682 -1034 2154 -975
rect 2097 -1359 2154 -1034
<< metal3 >>
rect 0 15633 348 17033
rect 257 11540 3861 11699
rect 3845 9433 4055 11339
rect 222 3781 1617 3843
rect 3938 2529 4055 3483
rect 3945 444 4055 762
use din_512x8m81  din_512x8m81_0
timestamp 1763476864
transform 1 0 226 0 1 5803
box -156 -50 1824 6415
use M2_M1$$45012012_512x8m81  M2_M1$$45012012_512x8m81_0
timestamp 1763476864
transform 1 0 1789 0 1 11647
box -562 -46 562 46
use M2_M1$$45013036_512x8m81  M2_M1$$45013036_512x8m81_0
timestamp 1763476864
transform 1 0 2870 0 1 11647
box -266 -46 266 46
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_0
timestamp 1763476864
transform 0 -1 3614 1 0 4199
box -63 -34 63 34
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_1
timestamp 1763476864
transform 0 -1 3273 1 0 4199
box -63 -34 63 34
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_2
timestamp 1763476864
transform 1 0 669 0 1 252
box -63 -34 63 34
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_0
timestamp 1763476864
transform 1 0 2126 0 1 -1300
box -34 -63 34 63
use m2_saout01_512x8m81  m2_saout01_512x8m81_0
timestamp 1763476864
transform 1 0 480 0 1 20286
box -102 -44 3491 1507
use M3_M2$$43370540_512x8m81  M3_M2$$43370540_512x8m81_0
timestamp 1763476864
transform 1 0 2870 0 1 11647
box -266 -46 266 46
use M3_M2$$44741676_512x8m81  M3_M2$$44741676_512x8m81_0
timestamp 1763476864
transform 1 0 1759 0 1 11647
box -562 -46 562 46
use M3_M2431059130207_512x8m81  M3_M2431059130207_512x8m81_0
timestamp 1763476864
transform 1 0 1554 0 1 3812
box -63 -35 63 35
use mux821_512x8m81  mux821_512x8m81_0
timestamp 1763486358
transform 1 0 387 0 1 12003
box -575 93 4956 8484
use outbuf_oe_512x8m81  outbuf_oe_512x8m81_0
timestamp 1763476864
transform 1 0 442 0 1 4196
box -372 -251 3623 2326
use sa_512x8m81  sa_512x8m81_0
timestamp 1763476864
transform 1 0 442 0 1 6365
box -249 -137 3523 5747
use sacntl_2_512x8m81  sacntl_2_512x8m81_0
timestamp 1763476864
transform 1 0 442 0 1 356
box -371 -16 3623 3958
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_0
timestamp 1763476864
transform 1 0 1451 0 1 8980
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_1
timestamp 1763476864
transform 1 0 1451 0 1 8438
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_2
timestamp 1763476864
transform 1 0 1451 0 1 7797
box -9 0 73 215
use via1_R90_512x8m81  via1_R90_512x8m81_0
timestamp 1763476864
transform -1 0 3930 0 1 13423
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_1
timestamp 1763476864
transform 0 -1 439 1 0 11451
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_2
timestamp 1763476864
transform 0 -1 258 1 0 18907
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_3
timestamp 1763476864
transform -1 0 495 0 -1 13539
box 0 0 65 89
use via1_x2_512x8m81  via1_x2_512x8m81_0
timestamp 1763476864
transform -1 0 1644 0 -1 11518
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_1
timestamp 1763476864
transform -1 0 1103 0 -1 5011
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_2
timestamp 1763476864
transform 1 0 1579 0 1 2668
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_3
timestamp 1763476864
transform 1 0 3741 0 1 7312
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_4
timestamp 1763476864
transform 1 0 322 0 1 6111
box -8 0 72 222
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 3592 1 0 11775
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_1
timestamp 1763476864
transform 0 -1 1377 1 0 13448
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_2
timestamp 1763476864
transform 0 -1 2275 1 0 13454
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_3
timestamp 1763476864
transform 0 -1 3179 1 0 13454
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_4
timestamp 1763476864
transform 0 -1 647 1 0 6493
box -8 0 72 215
use via2_512x8m81  via2_512x8m81_0
timestamp 1763476864
transform -1 0 619 0 1 13417
box 0 0 65 92
use via2_512x8m81  via2_512x8m81_1
timestamp 1763476864
transform -1 0 1207 0 1 13667
box 0 0 65 92
use via2_512x8m81  via2_512x8m81_2
timestamp 1763476864
transform -1 0 1396 0 1 13896
box 0 0 65 92
use via2_512x8m81  via2_512x8m81_3
timestamp 1763476864
transform -1 0 3011 0 1 14925
box 0 0 65 92
use via2_512x8m81  via2_512x8m81_4
timestamp 1763476864
transform -1 0 3200 0 1 15166
box 0 0 65 92
use via2_512x8m81  via2_512x8m81_5
timestamp 1763476864
transform -1 0 3948 0 1 15409
box 0 0 65 92
use via2_512x8m81  via2_512x8m81_6
timestamp 1763476864
transform 1 0 2044 0 1 14154
box 0 0 65 92
use via2_512x8m81  via2_512x8m81_7
timestamp 1763476864
transform 1 0 2229 0 1 14696
box 0 0 65 92
use via2_x2_512x8m81  via2_x2_512x8m81_0
timestamp 1763476864
transform 1 0 271 0 1 16282
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_1
timestamp 1763476864
transform 1 0 26 0 1 16282
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_2
timestamp 1763476864
transform 1 0 1709 0 1 8980
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_3
timestamp 1763476864
transform 1 0 1709 0 1 8438
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_4
timestamp 1763476864
transform 1 0 1709 0 1 7797
box -9 0 74 222
use wen_wm1_512x8m81  wen_wm1_512x8m81_0
timestamp 1763486358
transform 1 0 225 0 1 -2023
box -133 -24 3461 2300
<< labels >>
rlabel metal3 s 653 20226 653 20226 4 vdd
port 10 nsew
rlabel metal2 s 3850 20107 3850 20107 4 b[7]
port 15 nsew
rlabel metal2 s 3124 20107 3124 20107 4 b[6]
port 16 nsew
rlabel metal2 s 2979 20107 2979 20107 4 b[5]
port 17 nsew
rlabel metal2 s 2259 20107 2259 20107 4 b[4]
port 18 nsew
rlabel metal2 s 2116 20107 2116 20107 4 b[3]
port 19 nsew
rlabel metal2 s 1388 20107 1388 20107 4 b[2]
port 20 nsew
rlabel metal2 s 1246 20107 1246 20107 4 b[1]
port 21 nsew
rlabel metal2 s 515 20108 515 20108 4 b[0]
port 22 nsew
rlabel metal2 s 3416 20108 3416 20108 4 bb[6]
port 23 nsew
rlabel metal2 s 3557 20113 3557 20113 4 bb[7]
port 24 nsew
rlabel metal2 s 2688 20108 2688 20108 4 bb[5]
port 25 nsew
rlabel metal2 s 2548 20108 2548 20108 4 bb[4]
port 27 nsew
rlabel metal2 s 1822 20113 1822 20113 4 bb[3]
port 28 nsew
rlabel metal2 s 1683 20111 1683 20111 4 bb[2]
port 29 nsew
rlabel metal2 s 813 20107 813 20107 4 bb[0]
port 30 nsew
rlabel metal2 s 957 20107 957 20107 4 bb[1]
port 31 nsew
rlabel metal3 s 616 1362 616 1362 4 men
port 8 nsew
rlabel metal3 s 261 1100 261 1100 4 vss
port 9 nsew
rlabel metal3 s 308 1865 308 1865 4 vss
port 9 nsew
rlabel metal3 s 567 14477 567 14477 4 ypass[4]
port 4 nsew
rlabel metal3 s 381 3030 381 3030 4 vdd
port 10 nsew
rlabel metal3 s 275 619 275 619 4 vdd
port 10 nsew
rlabel metal3 s 317 4648 317 4648 4 vss
port 9 nsew
rlabel metal3 s 307 8060 307 8060 4 vss
port 9 nsew
rlabel metal3 s 567 15149 567 15149 4 ypass[7]
port 7 nsew
rlabel metal3 s 567 14926 567 14926 4 ypass[6]
port 6 nsew
rlabel metal3 s 567 14704 567 14704 4 ypass[5]
port 5 nsew
rlabel metal3 s 567 14019 567 14019 4 ypass[3]
port 3 nsew
rlabel metal3 s 567 13796 567 13796 4 ypass[2]
port 2 nsew
rlabel metal3 s 567 13574 567 13574 4 ypass[1]
port 1 nsew
rlabel metal3 s 278 1360 278 1360 4 men
port 8 nsew
rlabel metal3 s 664 15745 664 15745 4 vss
port 9 nsew
rlabel metal3 s 333 12356 333 12356 4 vss
port 9 nsew
rlabel metal3 s 326 9974 326 9974 4 vdd
port 10 nsew
rlabel metal3 s 280 6448 280 6448 4 vdd
port 10 nsew
rlabel metal3 s 234 5497 234 5497 4 vdd
port 10 nsew
rlabel metal3 s 567 13349 567 13349 4 ypass[0]
port 11 nsew
flabel metal3 s 450 3811 450 3811 0 FreeSans 420 0 0 0 GWE
port 12 nsew
rlabel metal3 s 275 -74 275 -74 4 vdd
port 10 nsew
rlabel metal3 s 261 -893 261 -893 4 vss
port 9 nsew
rlabel metal3 s 261 -1291 261 -1291 4 vss
port 9 nsew
rlabel metal3 s 275 -1757 275 -1757 4 vdd
port 10 nsew
rlabel metal3 s 261 -622 261 -622 4 vss
port 9 nsew
flabel metal3 s 493 -1063 493 -1063 0 FreeSans 420 0 0 0 GWEN
port 13 nsew
rlabel metal1 s 695 19292 695 19292 4 pcb
port 32 nsew
rlabel metal1 s 488 6159 488 6159 4 datain
port 14 nsew
rlabel metal1 s 695 19291 695 19291 4 pcb
port 32 nsew
rlabel metal1 s 653 13049 653 13049 4 vdd
port 10 nsew
flabel metal1 s 496 -2000 496 -2000 0 FreeSans 420 0 0 0 WEN
port 33 nsew
rlabel metal2 s 965 1150 965 1150 4 q
port 26 nsew
rlabel metal2 s 965 1126 965 1126 4 q
port 26 nsew
rlabel metal2 s 352 1477 352 1477 4 datain
port 14 nsew
<< properties >>
string path 10.130 4.930 10.130 -9.675 15.190 -9.675 15.190 -12.125 
<< end >>
