magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -70 280 70 287
rect -70 -280 -63 280
rect 63 -280 70 280
rect -70 -287 70 -280
<< via2 >>
rect -63 -280 63 280
<< metal3 >>
rect -70 280 70 287
rect -70 -280 -63 280
rect 63 -280 70 280
rect -70 -287 70 -280
<< end >>
