magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -113 627 113 634
rect -113 -627 -106 627
rect 106 -627 113 627
rect -113 -634 113 -627
<< via2 >>
rect -106 -627 106 627
<< metal3 >>
rect -113 627 113 634
rect -113 -627 -106 627
rect 106 -627 113 627
rect -113 -634 113 -627
<< end >>
