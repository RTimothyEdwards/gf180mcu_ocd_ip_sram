magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal1 >>
rect -330 105 330 113
rect -330 -105 -322 105
rect 322 -105 330 105
rect -330 -113 330 -105
<< via1 >>
rect -322 -105 322 105
<< metal2 >>
rect -330 105 330 113
rect -330 -105 -322 105
rect 322 -105 330 105
rect -330 -113 330 -105
<< end >>
