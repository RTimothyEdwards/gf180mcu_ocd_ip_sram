magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< nwell >>
rect -426 -86 1422 526
<< pmos >>
rect -252 0 -196 440
rect -92 0 -36 440
rect 69 0 125 440
rect 229 0 285 440
rect 390 0 446 440
rect 550 0 606 440
rect 711 0 767 440
rect 871 0 927 440
rect 1032 0 1088 440
rect 1192 0 1248 440
<< pdiff >>
rect -340 427 -252 440
rect -340 13 -327 427
rect -281 13 -252 427
rect -340 0 -252 13
rect -196 427 -92 440
rect -196 13 -167 427
rect -121 13 -92 427
rect -196 0 -92 13
rect -36 427 69 440
rect -36 13 -7 427
rect 39 13 69 427
rect -36 0 69 13
rect 125 427 229 440
rect 125 13 154 427
rect 200 13 229 427
rect 125 0 229 13
rect 285 427 390 440
rect 285 13 314 427
rect 360 13 390 427
rect 285 0 390 13
rect 446 427 550 440
rect 446 13 475 427
rect 521 13 550 427
rect 446 0 550 13
rect 606 427 711 440
rect 606 13 635 427
rect 681 13 711 427
rect 606 0 711 13
rect 767 427 871 440
rect 767 13 796 427
rect 842 13 871 427
rect 767 0 871 13
rect 927 427 1032 440
rect 927 13 956 427
rect 1002 13 1032 427
rect 927 0 1032 13
rect 1088 427 1192 440
rect 1088 13 1117 427
rect 1163 13 1192 427
rect 1088 0 1192 13
rect 1248 427 1336 440
rect 1248 13 1277 427
rect 1323 13 1336 427
rect 1248 0 1336 13
<< pdiffc >>
rect -327 13 -281 427
rect -167 13 -121 427
rect -7 13 39 427
rect 154 13 200 427
rect 314 13 360 427
rect 475 13 521 427
rect 635 13 681 427
rect 796 13 842 427
rect 956 13 1002 427
rect 1117 13 1163 427
rect 1277 13 1323 427
<< polysilicon >>
rect -252 440 -196 484
rect -92 440 -36 484
rect 69 440 125 484
rect 229 440 285 484
rect 390 440 446 484
rect 550 440 606 484
rect 711 440 767 484
rect 871 440 927 484
rect 1032 440 1088 484
rect 1192 440 1248 484
rect -252 -44 -196 0
rect -92 -44 -36 0
rect 69 -44 125 0
rect 229 -44 285 0
rect 390 -44 446 0
rect 550 -44 606 0
rect 711 -44 767 0
rect 871 -44 927 0
rect 1032 -44 1088 0
rect 1192 -44 1248 0
<< metal1 >>
rect -327 427 -281 440
rect -327 0 -281 13
rect -167 427 -121 440
rect -167 0 -121 13
rect -7 427 39 440
rect -7 0 39 13
rect 154 427 200 440
rect 154 0 200 13
rect 314 427 360 440
rect 314 0 360 13
rect 475 427 521 440
rect 475 0 521 13
rect 635 427 681 440
rect 635 0 681 13
rect 796 427 842 440
rect 796 0 842 13
rect 956 427 1002 440
rect 956 0 1002 13
rect 1117 427 1163 440
rect 1117 0 1163 13
rect 1277 427 1323 440
rect 1277 0 1323 13
<< labels >>
flabel pdiffc 498 220 498 220 0 FreeSans 186 0 0 0 D
flabel pdiffc -292 220 -292 220 0 FreeSans 186 0 0 0 S
flabel pdiffc -132 220 -132 220 0 FreeSans 186 0 0 0 D
flabel pdiffc 28 220 28 220 0 FreeSans 186 0 0 0 S
flabel pdiffc 189 220 189 220 0 FreeSans 186 0 0 0 D
flabel pdiffc 349 220 349 220 0 FreeSans 186 0 0 0 S
flabel pdiffc 646 220 646 220 0 FreeSans 186 0 0 0 S
flabel pdiffc 807 220 807 220 0 FreeSans 186 0 0 0 D
flabel pdiffc 1128 220 1128 220 0 FreeSans 186 0 0 0 D
flabel pdiffc 967 220 967 220 0 FreeSans 186 0 0 0 S
flabel pdiffc 1288 220 1288 220 0 FreeSans 186 0 0 0 S
<< end >>
