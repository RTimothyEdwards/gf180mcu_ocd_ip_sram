magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect 407 -103 2148 777
rect 3304 -49 5064 754
rect 5922 -64 6342 789
rect 9980 -49 13719 758
rect 14873 -2 16844 750
rect 16534 -103 16844 -2
<< nmos >>
rect 9450 501 9744 557
rect 2520 190 2986 246
rect 9450 366 9744 422
rect 9450 224 9744 280
rect 14035 190 14501 246
<< ndiff >>
rect 9450 641 9744 678
rect 9450 595 9474 641
rect 9721 595 9744 641
rect 9450 557 9744 595
rect 9450 422 9744 501
rect 2520 281 2986 345
rect 2520 246 2986 270
rect 2520 161 2986 190
rect 2520 115 2535 161
rect 2969 115 2986 161
rect 9450 280 9744 366
rect 9450 186 9744 224
rect 9450 140 9474 186
rect 9721 140 9744 186
rect 14035 246 14501 345
rect 14035 161 14501 190
rect 9450 123 9744 140
rect 2520 102 2986 115
rect 14035 115 14071 161
rect 14481 115 14501 161
rect 14035 98 14501 115
<< ndiffc >>
rect 9474 595 9721 641
rect 2535 115 2969 161
rect 9474 140 9721 186
rect 14071 115 14481 161
<< nsubdiff >>
rect 10612 678 12713 686
rect 507 566 616 673
rect 4160 570 4519 667
rect 507 63 538 566
rect 584 63 616 566
rect 10612 590 12853 678
rect 10612 492 10643 590
rect 12681 581 12853 590
rect 12681 492 12713 581
rect 16634 566 16744 673
rect 10612 459 12713 492
rect 507 0 616 63
rect 16634 63 16666 566
rect 16712 63 16744 566
rect 16634 0 16744 63
<< nsubdiffcont >>
rect 538 63 584 566
rect 10643 492 12681 590
rect 16666 63 16712 566
<< polysilicon >>
rect 2186 510 2479 566
rect 6854 534 6966 566
rect 9797 557 10032 565
rect 6853 527 6966 534
rect 6854 510 6966 527
rect 9065 501 9450 557
rect 9744 509 10032 557
rect 9744 501 9846 509
rect 9065 492 9189 501
rect 14545 510 14925 566
rect 2186 350 2479 406
rect 3310 304 3618 360
rect 3310 246 3351 304
rect 2476 190 2520 246
rect 2986 200 3351 246
rect 2986 190 3618 200
rect 3310 144 3618 190
rect 4218 135 4295 375
rect 4391 360 4458 375
rect 4391 304 4617 360
rect 5749 317 5831 373
rect 9401 366 9450 422
rect 9744 406 9828 422
rect 9744 366 10034 406
rect 4391 200 4458 304
rect 5756 213 5831 317
rect 9818 350 10034 366
rect 9401 224 9450 280
rect 9744 246 9886 280
rect 9744 224 10034 246
rect 4391 144 4617 200
rect 5749 157 5831 213
rect 6286 150 6426 206
rect 6571 150 6591 206
rect 9820 190 10034 224
rect 10362 190 10466 246
rect 12739 144 12810 375
rect 13407 304 13710 360
rect 14545 350 14797 406
rect 14869 349 14925 405
rect 13669 246 13710 304
rect 13669 200 14035 246
rect 13407 190 14035 200
rect 14501 190 14545 246
rect 13407 144 13710 190
rect 14869 189 14925 245
<< metal1 >>
rect 470 566 675 676
rect 4140 576 4587 660
rect 5279 583 5544 676
rect 16576 672 16781 676
rect 470 63 538 566
rect 584 347 675 566
rect 584 264 1290 347
rect 584 63 675 264
rect 2137 177 2184 434
rect 4223 378 4696 462
rect 4924 378 5268 462
rect 3192 217 4169 302
rect 2523 177 2985 178
rect 3192 177 3274 217
rect 2137 161 3274 177
rect 2137 115 2535 161
rect 2969 115 3274 161
rect 2137 113 3274 115
rect 4223 138 4305 378
rect 4365 194 4458 322
rect 4924 217 5426 300
rect 470 -46 675 63
rect 4223 54 4701 138
rect 4924 54 5268 138
rect 5777 124 5825 315
rect 6027 217 6243 672
rect 6361 588 7488 672
rect 9457 655 9739 672
rect 8321 641 9739 655
rect 8321 604 9474 641
rect 9457 595 9474 604
rect 9721 595 9739 641
rect 6361 285 6442 588
rect 9457 585 9739 595
rect 10435 590 12928 672
rect 10435 588 10643 590
rect 6617 435 6630 481
rect 6361 239 6464 285
rect 6663 209 6776 359
rect 6583 186 6776 209
rect 6889 186 6970 513
rect 7219 416 9184 510
rect 10626 492 10643 588
rect 12681 588 12928 590
rect 16435 588 16781 672
rect 12681 492 12699 588
rect 16576 566 16781 588
rect 10626 473 12699 492
rect 9940 425 10126 472
rect 9775 347 9893 418
rect 8277 254 9893 347
rect 9940 186 10021 425
rect 6583 140 9474 186
rect 9721 140 10159 186
rect 10497 178 12582 272
rect 13332 217 13829 300
rect 3126 -26 3234 51
rect 5777 40 6523 124
rect 6583 102 10159 140
rect 13748 177 13829 217
rect 14803 177 14863 517
rect 16576 347 16666 566
rect 15739 264 16666 347
rect 13748 161 14863 177
rect 13748 115 14071 161
rect 14481 115 14863 161
rect 13748 112 14863 115
rect 16576 63 16666 264
rect 16712 63 16781 566
rect 13786 -20 13895 51
rect 16576 -46 16781 63
<< metal2 >>
rect 486 -70 1739 681
rect 1830 113 2046 520
rect 2328 261 2580 535
rect 2676 -70 3234 735
rect 3308 -70 4207 735
rect 4365 207 4455 359
rect 4522 -70 5138 735
rect 5213 48 5429 473
rect 5505 -70 5922 735
rect 5994 -70 6450 735
rect 6532 147 6622 510
rect 6867 -70 7084 735
rect 7219 -156 7374 735
rect 7483 -156 7639 735
rect 7748 -156 7903 744
rect 8012 -156 8167 744
rect 8277 -156 8432 744
rect 8541 -156 8696 744
rect 8806 -156 8960 744
rect 9070 -156 9225 744
rect 9310 -143 9911 735
rect 10047 -143 10486 735
rect 10577 -156 10731 744
rect 10840 -156 10996 744
rect 11105 -156 11260 744
rect 11370 -156 11524 744
rect 11634 -156 11789 744
rect 11898 -156 12054 744
rect 12163 -156 12318 744
rect 12427 -156 12582 744
rect 12870 -70 13710 735
rect 13786 -70 14356 735
rect 14441 251 14658 520
rect 14974 98 15191 515
rect 15276 -70 16765 735
<< metal3 >>
rect 230 547 16952 688
rect 230 251 2580 392
rect 4370 308 6745 402
rect 14441 251 16952 392
rect 5213 147 12798 240
rect 230 -58 16952 82
use M1_NWELL07_512x8m81  M1_NWELL07_512x8m81_0
timestamp 1763476864
transform 1 0 6132 0 1 618
box -210 -159 210 159
use M1_NWELL4310591302032_512x8m81  M1_NWELL4310591302032_512x8m81_0
timestamp 1763476864
transform 1 0 4341 0 1 618
box -126 -85 127 87
use M1_PACTIVE03_512x8m81  M1_PACTIVE03_512x8m81_0
timestamp 1763476864
transform 1 0 3174 0 -1 12
box -54 -56 54 56
use M1_PACTIVE43105913020106_51_0  M1_PACTIVE43105913020106_51_0_0
timestamp 1763476864
transform 1 0 5467 0 1 618
box -193 -36 193 36
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_0
timestamp 1763476864
transform 0 1 10591 -1 0 233
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_1
timestamp 1763476864
transform 1 0 4421 0 1 257
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_2
timestamp 1763476864
transform 1 0 5801 0 1 259
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_3
timestamp 1763476864
transform 1 0 12768 0 1 276
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_4
timestamp 1763476864
transform 1 0 4265 0 1 257
box -36 -126 60 122
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1763476864
transform 1 0 6930 0 1 474
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1763476864
transform 1 0 6624 0 1 179
box -36 -36 36 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_0
timestamp 1763476864
transform 1 0 9836 0 1 394
box -62 -36 62 36
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_1
timestamp 1763476864
transform 1 0 9127 0 1 501
box -62 -36 62 36
use M1_POLY243105913020105_512x8m81  M1_POLY243105913020105_512x8m81_0
timestamp 1763476864
transform 1 0 14833 0 1 350
box -36 -161 36 161
use M1_POLY243105913020105_512x8m81  M1_POLY243105913020105_512x8m81_1
timestamp 1763476864
transform 1 0 2154 0 1 388
box -36 -161 36 161
use M1_PSUB$$45111340_512x8m81  M1_PSUB$$45111340_512x8m81_0
timestamp 1763476864
transform -1 0 13845 0 -1 12
box -56 -58 56 58
use M1_PSUB_05_512x8m81  M1_PSUB_05_512x8m81_0
timestamp 1763476864
transform 1 0 8038 0 1 618
box -775 -58 775 58
use M2_M1$$45004844_512x8m81  M2_M1$$45004844_512x8m81_0
timestamp 1763476864
transform 1 0 14125 0 1 618
box -193 -46 193 46
use M2_M1$$46894124_512x8m81  M2_M1$$46894124_512x8m81_0
timestamp 1763476864
transform 1 0 4410 0 1 254
box -44 -46 45 46
use M2_M1$$201262124_512x8m81  M2_M1$$201262124_512x8m81_0
timestamp 1763476864
transform 1 0 10266 0 1 291
box -119 -46 119 46
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_0
timestamp 1763476864
transform 1 0 4410 0 1 254
box -44 -46 44 46
use M2_M1$$202394668_512x8m81  M2_M1$$202394668_512x8m81_1
timestamp 1763476864
transform 1 0 6577 0 1 463
box -44 -46 44 46
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_0
timestamp 1763476864
transform 1 0 12752 0 1 269
box -45 -122 45 123
use M2_M1$$204402732_512x8m81  M2_M1$$204402732_512x8m81_0
timestamp 1763476864
transform 1 0 16020 0 -1 12
box -709 -46 709 46
use M2_M1$$204402732_512x8m81  M2_M1$$204402732_512x8m81_1
timestamp 1763476864
transform 1 0 16020 0 1 618
box -709 -46 709 46
use M2_M1$$204402732_512x8m81  M2_M1$$204402732_512x8m81_2
timestamp 1763476864
transform 1 0 997 0 1 12
box -709 -46 709 46
use M2_M1$$204402732_512x8m81  M2_M1$$204402732_512x8m81_3
timestamp 1763476864
transform 1 0 997 0 1 618
box -709 -46 709 46
use M2_M1$$204403756_512x8m81  M2_M1$$204403756_512x8m81_0
timestamp 1763476864
transform 1 0 5322 0 1 427
box -107 -46 107 46
use M2_M1$$204403756_512x8m81  M2_M1$$204403756_512x8m81_1
timestamp 1763476864
transform 1 0 6975 0 1 618
box -107 -46 107 46
use M2_M1$$204403756_512x8m81  M2_M1$$204403756_512x8m81_2
timestamp 1763476864
transform 1 0 15082 0 1 468
box -107 -46 107 46
use M2_M1$$204403756_512x8m81  M2_M1$$204403756_512x8m81_3
timestamp 1763476864
transform 1 0 13895 0 -1 12
box -107 -46 107 46
use M2_M1$$204403756_512x8m81  M2_M1$$204403756_512x8m81_4
timestamp 1763476864
transform 1 0 6134 0 1 618
box -107 -46 107 46
use M2_M1$$204403756_512x8m81  M2_M1$$204403756_512x8m81_5
timestamp 1763476864
transform 1 0 3126 0 -1 12
box -107 -46 107 46
use M2_M1$$204403756_512x8m81  M2_M1$$204403756_512x8m81_6
timestamp 1763476864
transform 1 0 5322 0 1 95
box -107 -46 107 46
use M2_M1$$204403756_512x8m81  M2_M1$$204403756_512x8m81_7
timestamp 1763476864
transform 1 0 14549 0 1 473
box -107 -46 107 46
use M2_M1$$204403756_512x8m81  M2_M1$$204403756_512x8m81_8
timestamp 1763476864
transform 1 0 1938 0 1 471
box -107 -46 107 46
use M2_M1$$204403756_512x8m81  M2_M1$$204403756_512x8m81_9
timestamp 1763476864
transform 1 0 1938 0 1 151
box -107 -46 107 46
use M2_M1$$204403756_512x8m81  M2_M1$$204403756_512x8m81_10
timestamp 1763476864
transform 1 0 2471 0 1 493
box -107 -46 107 46
use M2_M1$$204403756_512x8m81  M2_M1$$204403756_512x8m81_11
timestamp 1763476864
transform 1 0 15082 0 1 144
box -107 -46 107 46
use M2_M1$$204404780_512x8m81  M2_M1$$204404780_512x8m81_0
timestamp 1763476864
transform 1 0 9610 0 1 618
box -266 -46 266 46
use M2_M1$$204404780_512x8m81  M2_M1$$204404780_512x8m81_1
timestamp 1763476864
transform 1 0 2956 0 1 618
box -266 -46 266 46
use M2_M1$$204404780_512x8m81  M2_M1$$204404780_512x8m81_2
timestamp 1763476864
transform 1 0 4830 0 1 259
box -266 -46 266 46
use M2_M1$$204405804_512x8m81  M2_M1$$204405804_512x8m81_0
timestamp 1763476864
transform 1 0 2848 0 1 306
box -171 -46 171 46
use M2_M1$$204406828_512x8m81  M2_M1$$204406828_512x8m81_0
timestamp 1763476864
transform 1 0 13290 0 1 618
box -414 -46 414 46
use M2_M1$$204406828_512x8m81  M2_M1$$204406828_512x8m81_1
timestamp 1763476864
transform 1 0 3758 0 1 618
box -414 -46 414 46
use M2_M1$$204407852_512x8m81  M2_M1$$204407852_512x8m81_0
timestamp 1763476864
transform 1 0 3763 0 1 418
box -340 -46 340 46
use M2_M1$$204407852_512x8m81  M2_M1$$204407852_512x8m81_1
timestamp 1763476864
transform 1 0 3763 0 1 96
box -340 -46 340 46
use M2_M1$$204407852_512x8m81  M2_M1$$204407852_512x8m81_2
timestamp 1763476864
transform 1 0 13290 0 1 420
box -340 -46 340 46
use M2_M1$$204407852_512x8m81  M2_M1$$204407852_512x8m81_3
timestamp 1763476864
transform 1 0 13290 0 1 96
box -340 -46 340 46
use M2_M1$$204408876_512x8m81  M2_M1$$204408876_512x8m81_0
timestamp 1763476864
transform 1 0 10266 0 1 618
box -193 -46 193 46
use M2_M1$$204408876_512x8m81  M2_M1$$204408876_512x8m81_1
timestamp 1763476864
transform 1 0 14093 0 1 306
box -193 -46 193 46
use M2_M1$$204408876_512x8m81  M2_M1$$204408876_512x8m81_2
timestamp 1763476864
transform 1 0 5714 0 1 618
box -193 -46 193 46
use M2_M1$02_R270_512x8m81  M2_M1$02_R270_512x8m81_0
timestamp 1763476864
transform 0 -1 6731 1 0 247
box -112 -45 112 45
use M3_M2$$201251884_512x8m81  M3_M2$$201251884_512x8m81_0
timestamp 1763476864
transform 1 0 14071 0 -1 12
box -266 -46 266 46
use M3_M2$$201251884_512x8m81  M3_M2$$201251884_512x8m81_1
timestamp 1763476864
transform 1 0 9610 0 -1 12
box -266 -46 266 46
use M3_M2$$201251884_512x8m81  M3_M2$$201251884_512x8m81_2
timestamp 1763476864
transform 1 0 2956 0 -1 12
box -266 -46 266 46
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_0
timestamp 1763476864
transform 1 0 12752 0 1 269
box -45 -122 45 123
use M3_M2$$204147756_512x8m81  M3_M2$$204147756_512x8m81_0
timestamp 1763476864
transform 1 0 10266 0 1 618
box -193 -46 193 46
use M3_M2$$204147756_512x8m81  M3_M2$$204147756_512x8m81_1
timestamp 1763476864
transform 1 0 5714 0 -1 12
box -193 -46 193 46
use M3_M2$$204398636_512x8m81  M3_M2$$204398636_512x8m81_0
timestamp 1763476864
transform 1 0 6731 0 1 355
box -44 -46 45 46
use M3_M2$$204398636_512x8m81  M3_M2$$204398636_512x8m81_1
timestamp 1763476864
transform 1 0 4410 0 1 355
box -44 -46 45 46
use M3_M2$$204398636_512x8m81  M3_M2$$204398636_512x8m81_2
timestamp 1763476864
transform 1 0 6577 0 1 193
box -44 -46 45 46
use M3_M2$$204399660_512x8m81  M3_M2$$204399660_512x8m81_0
timestamp 1763476864
transform 1 0 16020 0 1 618
box -709 -46 709 46
use M3_M2$$204399660_512x8m81  M3_M2$$204399660_512x8m81_1
timestamp 1763476864
transform 1 0 997 0 1 618
box -709 -46 709 46
use M3_M2$$204400684_512x8m81  M3_M2$$204400684_512x8m81_0
timestamp 1763476864
transform 1 0 6975 0 -1 12
box -108 -46 108 46
use M3_M2$$204400684_512x8m81  M3_M2$$204400684_512x8m81_1
timestamp 1763476864
transform 1 0 5322 0 1 193
box -108 -46 108 46
use M3_M2$$204400684_512x8m81  M3_M2$$204400684_512x8m81_2
timestamp 1763476864
transform 1 0 1938 0 1 326
box -108 -46 108 46
use M3_M2$$204400684_512x8m81  M3_M2$$204400684_512x8m81_3
timestamp 1763476864
transform 1 0 2471 0 1 302
box -108 -46 108 46
use M3_M2$$204400684_512x8m81  M3_M2$$204400684_512x8m81_4
timestamp 1763476864
transform 1 0 14549 0 1 322
box -108 -46 108 46
use M3_M2$$204400684_512x8m81  M3_M2$$204400684_512x8m81_5
timestamp 1763476864
transform 1 0 6134 0 1 618
box -108 -46 108 46
use M3_M2$$204400684_512x8m81  M3_M2$$204400684_512x8m81_6
timestamp 1763476864
transform 1 0 15082 0 1 322
box -108 -46 108 46
use M3_M2$$204401708_512x8m81  M3_M2$$204401708_512x8m81_0
timestamp 1763476864
transform 1 0 13290 0 1 618
box -414 -46 414 46
use M3_M2$$204401708_512x8m81  M3_M2$$204401708_512x8m81_1
timestamp 1763476864
transform 1 0 3758 0 1 618
box -414 -46 414 46
use nmos_1p2_02_R270_512x8m81  nmos_1p2_02_R270_512x8m81_0
timestamp 1763476864
transform 0 -1 6834 1 0 524
box -102 -44 130 249
use nmos_5p043105913020106_512x8m81  nmos_5p043105913020106_512x8m81_0
timestamp 1763476864
transform 0 -1 6528 1 0 150
box -92 -44 148 105
use nmos_5p043105913020107_512x8m81  nmos_5p043105913020107_512x8m81_0
timestamp 1763476864
transform 0 -1 2986 -1 0 538
box -116 -44 276 510
use nmos_5p043105913020107_512x8m81  nmos_5p043105913020107_512x8m81_1
timestamp 1763476864
transform 0 1 14035 -1 0 538
box -116 -44 276 510
use nmos_5p043105913020109_512x8m81  nmos_5p043105913020109_512x8m81_0
timestamp 1763476864
transform 0 -1 5706 1 0 185
box -116 -44 276 352
use pmos_1p2_01_R270_512x8m81  pmos_1p2_01_R270_512x8m81_0
timestamp 1763476864
transform 0 1 12852 1 0 186
box -246 -93 428 606
use pmos_1p2_01_R270_512x8m81  pmos_1p2_01_R270_512x8m81_1
timestamp 1763476864
transform 0 -1 4174 1 0 186
box -246 -93 428 606
use pmos_1p2_02_R270_512x8m81  pmos_1p2_02_R270_512x8m81_0
timestamp 1763476864
transform 0 -1 4967 1 0 186
box -216 -86 398 394
use pmos_1p2_03_R270_512x8m81  pmos_1p2_03_R270_512x8m81_0
timestamp 1763476864
transform 0 -1 2052 1 0 259
box -244 -138 481 1088
use pmos_5p043105913020103_512x8m81  pmos_5p043105913020103_512x8m81_0
timestamp 1763476864
transform 0 1 14969 1 0 245
box -230 -86 495 1019
use pmos_5p043105913020105_512x8m81  pmos_5p043105913020105_512x8m81_1
timestamp 1763476864
transform 0 1 10076 1 0 350
box -174 -86 230 330
use pmos_5p043105913020105_512x8m81  pmos_5p043105913020105_512x8m81_2
timestamp 1763476864
transform 0 1 10076 1 0 190
box -174 -86 230 330
use pmos_5p043105913020105_512x8m81  pmos_5p043105913020105_512x8m81_3
timestamp 1763476864
transform 0 1 10076 1 0 510
box -174 -86 230 330
use pmos_5p043105913020110_512x8m81  pmos_5p043105913020110_512x8m81_0
timestamp 1763476864
transform 0 -1 6245 1 0 150
box -174 -86 230 234
<< labels >>
rlabel metal3 s 16396 322 16396 322 4 RWL
port 3 nsew
rlabel metal2 s 4830 598 4830 598 4 men
port 5 nsew
rlabel metal1 s 9143 463 9143 463 4 xc
port 6 nsew
rlabel metal1 s 9143 301 9143 301 4 xb
port 7 nsew
rlabel metal1 s 10542 225 10542 225 4 xa
port 8 nsew
rlabel metal3 s 811 322 811 322 4 LWL
port 4 nsew
rlabel metal3 s 366 618 366 618 4 vdd
port 2 nsew
rlabel metal3 s 366 12 366 12 4 vss
port 1 nsew
rlabel metal3 s 366 36 366 36 2 vss
port 1 nsew
<< end >>
