magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nmos >>
rect 0 0 56 423
<< ndiff >>
rect -88 410 0 423
rect -88 13 -75 410
rect -29 13 0 410
rect -88 0 0 13
rect 56 410 144 423
rect 56 13 85 410
rect 131 13 144 410
rect 56 0 144 13
<< ndiffc >>
rect -75 13 -29 410
rect 85 13 131 410
<< polysilicon >>
rect 0 423 56 467
rect 0 -44 56 0
<< metal1 >>
rect -75 410 -29 423
rect -75 0 -29 13
rect 85 410 131 423
rect 85 0 131 13
<< labels >>
flabel ndiffc -40 211 -40 211 0 FreeSans 93 0 0 0 S
flabel ndiffc 96 211 96 211 0 FreeSans 93 0 0 0 D
<< end >>
