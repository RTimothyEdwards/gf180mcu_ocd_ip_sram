magic
tech gf180mcuD
magscale 1 10
timestamp 1764692000
<< nwell >>
rect 4608 38931 6692 39578
rect 9694 39386 10581 39589
rect 9694 39332 10808 39386
rect 7130 38937 7550 38988
rect 9695 38942 10808 39332
rect 4608 38896 6273 38931
rect 11564 38909 14760 39558
<< nsubdiff >>
rect 1486 39007 1594 39169
rect 17843 39021 17952 39169
rect 17842 38880 18051 39021
rect 17842 38794 18034 38880
<< polysilicon >>
rect 4589 39256 5251 39312
rect 4589 39180 4661 39256
rect 4485 39152 4661 39180
rect 7730 39172 7969 39180
rect 4485 39124 5251 39152
rect 7730 39124 8050 39172
rect 4592 39096 5251 39124
rect 7879 39116 8050 39124
rect 8358 39116 8451 39172
rect 9564 39137 9637 39435
rect 10754 39172 10826 39474
rect 12782 39256 13445 39312
rect 10713 39116 10826 39172
rect 10908 39117 11108 39172
rect 10908 39116 11028 39117
rect 11423 39116 11928 39173
rect 14707 39172 14779 39313
rect 12782 39096 13445 39152
rect 14707 39116 15356 39172
rect 14707 39096 14779 39116
<< metal1 >>
rect 1486 39067 2811 39462
rect 3026 39242 4435 39513
rect 4537 39162 5359 39246
rect 4537 39119 4618 39162
rect 1404 39007 2811 39067
rect 4368 39035 4618 39119
rect 6521 39119 6602 39335
rect 7969 39220 8339 39499
rect 9471 39405 9828 39499
rect 8404 39221 8919 39269
rect 9456 39221 10160 39269
rect 10687 39201 10961 39247
rect 11028 39197 11398 39499
rect 11659 39360 14659 39444
rect 11659 39231 12581 39360
rect 12788 39119 12849 39288
rect 14628 39181 14828 39228
rect 14926 39207 16342 39499
rect 6521 39035 8339 39119
rect 9499 39062 10170 39108
rect 11028 39035 12849 39119
rect 14746 39088 14828 39181
rect 14746 39042 15411 39088
rect 16625 39080 17952 39462
rect 16625 39007 18034 39080
rect 1404 38750 1506 39007
rect 17932 38793 18034 39007
<< metal2 >>
rect 1464 38795 2947 39539
rect 3885 38795 4442 39486
rect 4515 38795 5416 39486
rect 5730 38795 6346 39124
rect 6713 38795 7130 39486
rect 7193 38795 7658 39486
rect 8075 38795 8292 39486
rect 9795 39047 10181 39486
rect 8428 38757 8847 38900
rect 10518 38795 11120 39499
rect 14078 38795 14919 39486
rect 14994 38795 15565 39499
rect 16484 38795 17973 39539
rect 5992 -14 6083 78
rect 8988 -114 9079 -21
rect 9253 -114 9343 -21
rect 9517 -114 9608 -21
rect 9781 -114 9872 -21
rect 10046 -114 10136 -21
rect 10311 -114 10401 -21
rect 11817 -114 11907 -21
rect 12082 -114 12172 -21
rect 12345 -114 12436 -21
rect 12610 -114 12700 -21
rect 12875 -114 12965 -21
rect 13139 -114 13230 -21
rect 13403 -114 13493 -21
rect 13668 -114 13758 -21
<< metal3 >>
rect 48 39354 139 39447
rect 1443 39320 18161 39461
rect 428 39045 517 39138
rect 1443 39023 3714 39164
rect 5730 39031 9434 39124
rect 48 38754 139 38847
rect 9795 38808 9864 39068
rect 15655 39023 18161 39164
rect 18923 39045 19013 39138
rect 0 38452 89 38545
rect 19347 38452 19437 38545
rect 0 37834 89 37927
rect 19347 37834 19437 37927
rect 0 37240 89 37333
rect 19347 37240 19437 37333
rect 0 36621 89 36714
rect 19347 36622 19437 36715
rect 0 36028 89 36121
rect 19347 36028 19437 36121
rect 0 35410 89 35503
rect 19347 35410 19437 35503
rect 0 34816 89 34909
rect 19347 34816 19437 34909
rect 0 34198 89 34291
rect 19347 34198 19437 34291
rect 0 33604 89 33697
rect 19347 33604 19437 33697
rect 0 32986 89 33079
rect 19347 32986 19437 33079
rect 0 32393 89 32486
rect 19347 32392 19437 32485
rect 0 31774 89 31867
rect 19347 31774 19437 31867
rect 0 31181 89 31274
rect 19347 31180 19437 31273
rect 0 30562 89 30655
rect 19347 30562 19437 30655
rect 0 29969 89 30062
rect 19347 29969 19437 30062
rect 0 29350 89 29443
rect 19347 29351 19437 29444
rect 0 28756 89 28849
rect 19348 28756 19438 28849
rect 0 28138 89 28231
rect 19348 28139 19438 28232
rect 0 27544 89 27637
rect 19348 27545 19438 27638
rect 0 26926 89 27019
rect 19348 26926 19438 27019
rect 0 26333 89 26426
rect 19348 26332 19438 26425
rect 0 25714 89 25807
rect 19348 25714 19438 25807
rect 0 25119 89 25212
rect 19348 25120 19438 25213
rect 0 24502 89 24595
rect 19348 24502 19438 24595
rect 0 23908 89 24001
rect 19348 23908 19438 24001
rect 0 23289 89 23382
rect 19348 23290 19438 23383
rect 0 22696 89 22789
rect 19348 22696 19438 22789
rect 0 22077 89 22170
rect 19348 22077 19438 22170
rect 0 21484 89 21577
rect 19348 21484 19438 21577
rect 0 20865 89 20958
rect 19348 20866 19438 20959
rect 0 20273 89 20366
rect 19348 20272 19438 20365
rect 0 19653 89 19746
rect 19348 19652 19438 19745
rect 0 19059 89 19152
rect 19348 19059 19438 19152
rect 0 18441 89 18534
rect 19348 18443 19438 18536
rect 0 17847 89 17940
rect 19348 17847 19438 17940
rect 0 17231 89 17324
rect 19348 17231 19438 17324
rect 0 16631 89 16724
rect 19348 16635 19438 16728
rect 0 16015 89 16108
rect 19348 16019 19438 16112
rect 0 15423 89 15516
rect 19348 15423 19438 15516
rect 0 14807 89 14900
rect 19348 14807 19438 14900
rect 0 14211 89 14304
rect 19348 14211 19438 14304
rect 0 13595 89 13688
rect 19348 13595 19438 13688
rect 0 12999 89 13092
rect 19348 12999 19438 13092
rect 0 12383 89 12476
rect 19348 12383 19438 12476
rect 0 11787 89 11880
rect 19348 11787 19438 11880
rect 0 11171 89 11264
rect 19348 11171 19438 11264
rect 0 10575 89 10668
rect 19348 10575 19438 10668
rect 0 9959 89 10052
rect 19348 9959 19438 10052
rect 0 9363 89 9456
rect 19348 9363 19438 9456
rect 0 8747 89 8840
rect 19348 8747 19438 8840
rect 0 8150 89 8243
rect 19348 8151 19438 8244
rect 0 7534 89 7627
rect 19348 7535 19438 7628
rect 0 6939 89 7032
rect 19348 6939 19438 7032
rect 0 6323 89 6416
rect 19348 6323 19438 6416
rect 0 5727 89 5820
rect 19348 5727 19438 5820
rect 0 5111 89 5204
rect 19348 5111 19438 5204
rect 0 4515 89 4608
rect 19348 4515 19438 4608
rect 0 3899 89 3992
rect 19348 3899 19438 3992
rect 0 3301 89 3394
rect 19348 3301 19438 3394
rect 0 2685 89 2778
rect 19348 2685 19438 2778
rect 0 2091 89 2184
rect 19348 2091 19438 2184
rect 0 1475 89 1568
rect 19348 1475 19438 1568
rect 0 880 89 973
rect 19348 881 19438 974
rect 0 263 89 356
rect 19348 265 19438 358
use M1_NACTIVE_02_3v512x8m81  M1_NACTIVE_02_3v512x8m81_0
timestamp 1764525316
transform 1 0 9844 0 1 39457
box -54 -56 607 56
use M1_NWELL_01_3v512x8m81  M1_NWELL_01_3v512x8m81_0
timestamp 1764525316
transform 1 0 1540 0 1 39406
box -154 -501 1372 159
use M1_NWELL_01_3v512x8m81  M1_NWELL_01_3v512x8m81_1
timestamp 1764525316
transform -1 0 17897 0 1 39406
box -154 -501 1372 159
use M1_PACTIVE$10_3v512x8m81  M1_PACTIVE$10_3v512x8m81_0
timestamp 1764525316
transform 1 0 8024 0 1 39457
box -54 -56 1271 56
use M1_PACTIVE$10_3v512x8m81  M1_PACTIVE$10_3v512x8m81_1
timestamp 1764525316
transform 1 0 3073 0 1 39457
box -54 -56 1271 56
use M1_PACTIVE$10_3v512x8m81  M1_PACTIVE$10_3v512x8m81_2
timestamp 1764525316
transform 1 0 15032 0 1 39457
box -54 -56 1271 56
use M1_PACTIVE$11_3v512x8m81  M1_PACTIVE$11_3v512x8m81_0
timestamp 1764525316
transform 1 0 11102 0 1 39457
box -54 -56 275 56
use M1_POLY2$$204150828_3v512x8m81  M1_POLY2$$204150828_3v512x8m81_0
timestamp 1764525316
transform 1 0 6561 0 1 39204
box -46 -122 46 122
use M1_POLY24310591302019_3v512x8m81  M1_POLY24310591302019_3v512x8m81_0
timestamp 1764525316
transform 1 0 8428 0 1 39178
box -36 -80 36 78
use M1_POLY24310591302019_3v512x8m81  M1_POLY24310591302019_3v512x8m81_1
timestamp 1764525316
transform 0 -1 9598 1 0 39411
box -36 -80 36 78
use M1_POLY24310591302019_3v512x8m81  M1_POLY24310591302019_3v512x8m81_2
timestamp 1764525316
transform 1 0 10937 0 1 39206
box -36 -80 36 78
use M1_POLY24310591302019_3v512x8m81  M1_POLY24310591302019_3v512x8m81_3
timestamp 1764525316
transform 1 0 12819 0 1 39206
box -36 -80 36 78
use M1_POLY24310591302031_3v512x8m81  M1_POLY24310591302031_3v512x8m81_0
timestamp 1764525316
transform 1 0 10789 0 1 39444
box -36 -36 36 36
use M2_M1$$201262124_3v512x8m81  M2_M1$$201262124_3v512x8m81_0
timestamp 1764525316
transform 1 0 9590 0 1 39409
box -119 -46 119 46
use M2_M1$$204138540_3v512x8m81  M2_M1$$204138540_3v512x8m81_0
timestamp 1764525316
transform 1 0 7281 0 1 39239
box -45 -46 340 46
use M2_M1$$204138540_3v512x8m81  M2_M1$$204138540_3v512x8m81_1
timestamp 1764525316
transform 1 0 9841 0 1 39452
box -45 -46 340 46
use M2_M1$$204139564_3v512x8m81  M2_M1$$204139564_3v512x8m81_0
timestamp 1764525316
transform 1 0 8120 0 1 39419
box -45 -198 171 46
use M2_M1$$204140588_3v512x8m81  M2_M1$$204140588_3v512x8m81_0
timestamp 1764525316
transform 1 0 8651 0 1 39077
box -45 -46 783 46
use M2_M1$$204141612_3v512x8m81  M2_M1$$204141612_3v512x8m81_0
timestamp 1764525316
transform 1 0 10588 0 1 39452
box -45 -46 487 46
use M2_M1$$204141612_3v512x8m81  M2_M1$$204141612_3v512x8m81_1
timestamp 1764525316
transform 1 0 14123 0 1 39402
box -45 -46 487 46
use M2_M1$$204141612_3v512x8m81  M2_M1$$204141612_3v512x8m81_2
timestamp 1764525316
transform 1 0 14123 0 1 39077
box -45 -46 487 46
use M2_M1$$204220460_3v512x8m81  M2_M1$$204220460_3v512x8m81_0
timestamp 1764525316
transform 1 0 3079 0 1 39079
box -45 -46 635 46
use M2_M1$$204220460_3v512x8m81  M2_M1$$204220460_3v512x8m81_1
timestamp 1764525316
transform 1 0 4754 0 1 39367
box -45 -46 635 46
use M2_M1$$204220460_3v512x8m81  M2_M1$$204220460_3v512x8m81_2
timestamp 1764525316
transform 1 0 4754 0 1 39042
box -45 -46 635 46
use M2_M1$$204220460_3v512x8m81  M2_M1$$204220460_3v512x8m81_3
timestamp 1764525316
transform 1 0 15701 0 1 39077
box -45 -46 635 46
use M2_M1$$204221484_3v512x8m81  M2_M1$$204221484_3v512x8m81_0
timestamp 1764525316
transform 1 0 1509 0 1 39416
box -45 -351 1225 46
use M2_M1$$204221484_3v512x8m81  M2_M1$$204221484_3v512x8m81_1
timestamp 1764525316
transform -1 0 17928 0 1 39416
box -45 -351 1225 46
use M2_M1$$204222508_3v512x8m81  M2_M1$$204222508_3v512x8m81_0
timestamp 1764525316
transform 1 0 3947 0 1 39416
box -45 -198 487 46
use M2_M1$$204222508_3v512x8m81  M2_M1$$204222508_3v512x8m81_1
timestamp 1764525316
transform 1 0 15040 0 1 39416
box -45 -198 487 46
use M3_M2$$204142636_3v512x8m81  M3_M2$$204142636_3v512x8m81_0
timestamp 1764525316
transform 1 0 3947 0 1 39416
box -44 -46 487 46
use M3_M2$$204142636_3v512x8m81  M3_M2$$204142636_3v512x8m81_1
timestamp 1764525316
transform 1 0 5775 0 1 39077
box -44 -46 487 46
use M3_M2$$204142636_3v512x8m81  M3_M2$$204142636_3v512x8m81_2
timestamp 1764525316
transform 1 0 15040 0 1 39416
box -44 -46 487 46
use M3_M2$$204142636_3v512x8m81  M3_M2$$204142636_3v512x8m81_3
timestamp 1764525316
transform 1 0 15040 0 1 39416
box -44 -46 487 46
use M3_M2$$204143660_3v512x8m81  M3_M2$$204143660_3v512x8m81_0
timestamp 1764525316
transform 1 0 8120 0 1 39416
box -45 -46 171 46
use M3_M2$$204144684_3v512x8m81  M3_M2$$204144684_3v512x8m81_0
timestamp 1764525316
transform 1 0 3079 0 1 39079
box -45 -46 635 46
use M3_M2$$204144684_3v512x8m81  M3_M2$$204144684_3v512x8m81_1
timestamp 1764525316
transform 1 0 15701 0 1 39077
box -45 -46 635 46
use M3_M2$$204145708_3v512x8m81  M3_M2$$204145708_3v512x8m81_0
timestamp 1764525316
transform 1 0 8651 0 1 39077
box -45 -46 783 46
use M3_M2$$204146732_3v512x8m81  M3_M2$$204146732_3v512x8m81_0
timestamp 1764525316
transform 1 0 9841 0 1 39073
box -45 -46 340 46
use M3_M2$$204147756_3v512x8m81  M3_M2$$204147756_3v512x8m81_0
timestamp 1764525316
transform 1 0 8637 0 1 38786
box -193 -46 193 46
use nmos_1p2_01_R270_3v512x8m81  nmos_1p2_01_R270_3v512x8m81_0
timestamp 1764525316
transform 0 -1 9522 -1 0 39179
box -102 -44 130 659
use nmos_1p2_02_R90_3v512x8m81  nmos_1p2_02_R90_3v512x8m81_0
timestamp 1764525316
transform 0 -1 4442 1 0 39138
box -102 -44 130 987
use nmos_5p04310591302099_3v512x8m81  nmos_5p04310591302099_3v512x8m81_0
timestamp 1764525316
transform 0 -1 16342 1 0 39116
box -88 -44 144 987
use nmos_5p043105913020111_3v512x8m81  nmos_5p043105913020111_3v512x8m81_0
timestamp 1764525316
transform 0 -1 8339 1 0 39116
box -88 -44 144 291
use nmos_5p043105913020111_3v512x8m81  nmos_5p043105913020111_3v512x8m81_1
timestamp 1764525316
transform 0 -1 11398 1 0 39116
box -88 -44 144 291
use pmos_1p2_01_R90_3v512x8m81  pmos_1p2_01_R90_3v512x8m81_0
timestamp 1764525316
transform 0 -1 7702 1 0 39138
box -188 -86 216 701
use pmos_1p2_02_R90_3v512x8m81  pmos_1p2_02_R90_3v512x8m81_0
timestamp 1764525316
transform 0 -1 6471 1 0 39138
box -216 -86 348 1264
use pmos_1p2_02_R90_3v512x8m81  pmos_1p2_02_R90_3v512x8m81_1
timestamp 1764525316
transform 0 -1 14665 1 0 39138
box -216 -86 348 1264
use pmos_5p043105913020101_3v512x8m81  pmos_5p043105913020101_3v512x8m81_0
timestamp 1764525316
transform 0 -1 12581 1 0 39116
box -174 -86 230 701
use pmos_5p043105913020101_3v512x8m81  pmos_5p043105913020101_3v512x8m81_1
timestamp 1764525316
transform 0 -1 10712 1 0 39116
box -174 -86 230 701
use pmoscap_L1_W2_R270_3v512x8m81  pmoscap_L1_W2_R270_3v512x8m81_0
timestamp 1764692000
transform 0 -1 1542 -1 0 39446
box -88 -189 771 1517
use pmoscap_L1_W2_R270_3v512x8m81  pmoscap_L1_W2_R270_3v512x8m81_1
timestamp 1764692000
transform 0 1 17896 -1 0 39446
box -88 -189 771 1517
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_0
timestamp 1764525316
transform 0 1 17896 -1 0 10822
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_1
timestamp 1764525316
transform 0 1 17896 -1 0 9610
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_2
timestamp 1764525316
transform 0 1 17896 -1 0 8398
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_3
timestamp 1764525316
transform 0 1 17896 -1 0 7186
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_4
timestamp 1764525316
transform 0 1 17896 -1 0 5974
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_5
timestamp 1764525316
transform 0 1 17896 -1 0 4762
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_6
timestamp 1764525316
transform 0 1 17896 -1 0 3550
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_7
timestamp 1764525316
transform 0 1 17896 -1 0 2338
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_8
timestamp 1764525316
transform 0 1 17896 -1 0 1126
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_9
timestamp 1764525316
transform 0 1 17896 -1 0 19306
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_10
timestamp 1764525316
transform 0 1 17896 -1 0 18094
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_11
timestamp 1764525316
transform 0 1 17896 -1 0 16882
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_12
timestamp 1764525316
transform 0 1 17896 -1 0 15670
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_13
timestamp 1764525316
transform 0 1 17896 -1 0 14458
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_14
timestamp 1764525316
transform 0 1 17896 -1 0 13246
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_15
timestamp 1764525316
transform 0 1 17896 -1 0 12034
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_16
timestamp 1764525316
transform 0 -1 1542 -1 0 10822
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_17
timestamp 1764525316
transform 0 -1 1542 -1 0 9610
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_18
timestamp 1764525316
transform 0 -1 1542 -1 0 8398
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_19
timestamp 1764525316
transform 0 -1 1542 -1 0 7186
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_20
timestamp 1764525316
transform 0 -1 1542 -1 0 5974
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_21
timestamp 1764525316
transform 0 -1 1542 -1 0 4762
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_22
timestamp 1764525316
transform 0 -1 1542 -1 0 3550
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_23
timestamp 1764525316
transform 0 -1 1542 -1 0 2338
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_24
timestamp 1764525316
transform 0 -1 1542 -1 0 1126
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_25
timestamp 1764525316
transform 0 -1 1542 -1 0 19306
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_26
timestamp 1764525316
transform 0 -1 1542 -1 0 18094
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_27
timestamp 1764525316
transform 0 -1 1542 -1 0 16882
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_28
timestamp 1764525316
transform 0 -1 1542 -1 0 15670
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_29
timestamp 1764525316
transform 0 -1 1542 -1 0 14458
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_30
timestamp 1764525316
transform 0 -1 1542 -1 0 13246
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_31
timestamp 1764525316
transform 0 -1 1542 -1 0 12034
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_32
timestamp 1764525316
transform 0 -1 1542 -1 0 38698
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_33
timestamp 1764525316
transform 0 -1 1542 -1 0 37486
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_34
timestamp 1764525316
transform 0 -1 1542 -1 0 36274
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_35
timestamp 1764525316
transform 0 -1 1542 -1 0 35062
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_36
timestamp 1764525316
transform 0 -1 1542 -1 0 33850
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_37
timestamp 1764525316
transform 0 -1 1542 -1 0 32638
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_38
timestamp 1764525316
transform 0 -1 1542 -1 0 31426
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_39
timestamp 1764525316
transform 0 -1 1542 -1 0 30214
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_40
timestamp 1764525316
transform 0 -1 1542 -1 0 29002
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_41
timestamp 1764525316
transform 0 -1 1542 -1 0 27790
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_42
timestamp 1764525316
transform 0 -1 1542 -1 0 26578
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_43
timestamp 1764525316
transform 0 -1 1542 -1 0 25366
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_44
timestamp 1764525316
transform 0 -1 1542 -1 0 24154
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_45
timestamp 1764525316
transform 0 -1 1542 -1 0 22942
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_46
timestamp 1764525316
transform 0 -1 1542 -1 0 21730
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_47
timestamp 1764525316
transform 0 1 17896 -1 0 38698
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_48
timestamp 1764525316
transform 0 1 17896 -1 0 37486
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_49
timestamp 1764525316
transform 0 1 17896 -1 0 36274
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_50
timestamp 1764525316
transform 0 1 17896 -1 0 35062
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_51
timestamp 1764525316
transform 0 1 17896 -1 0 33850
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_52
timestamp 1764525316
transform 0 1 17896 -1 0 32638
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_53
timestamp 1764525316
transform 0 1 17896 -1 0 31426
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_54
timestamp 1764525316
transform 0 1 17896 -1 0 30214
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_55
timestamp 1764525316
transform 0 1 17896 -1 0 29002
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_56
timestamp 1764525316
transform 0 1 17896 -1 0 27790
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_57
timestamp 1764525316
transform 0 1 17896 -1 0 26578
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_58
timestamp 1764525316
transform 0 1 17896 -1 0 25366
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_59
timestamp 1764525316
transform 0 1 17896 -1 0 24154
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_60
timestamp 1764525316
transform 0 1 17896 -1 0 22942
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_61
timestamp 1764525316
transform 0 1 17896 -1 0 21730
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_62
timestamp 1764525316
transform 0 -1 1542 -1 0 20518
box -226 -219 1235 3808
use pmoscap_R270_3v512x8m81  pmoscap_R270_3v512x8m81_63
timestamp 1764525316
transform 0 1 17896 -1 0 20518
box -226 -219 1235 3808
use xdec32_3v512x8m81  xdec32_3v512x8m81_0
timestamp 1764692000
transform 1 0 1208 0 1 0
box 230 -159 16952 19575
use xdec32_468_3v512x8m81  xdec32_468_3v512x8m81_0
timestamp 1764692000
transform 1 0 1208 0 1 19392
box 230 -159 16952 19575
<< labels >>
rlabel metal2 s 10355 -67 10355 -67 4 xb[0]
port 133 nsew
rlabel metal2 s 10091 -67 10091 -67 4 xb[1]
port 134 nsew
rlabel metal2 s 9827 -67 9827 -67 4 xb[2]
port 135 nsew
rlabel metal2 s 9562 -67 9562 -67 4 xb[3]
port 136 nsew
rlabel metal2 s 11862 -67 11862 -67 4 xa[7]
port 137 nsew
rlabel metal2 s 12126 -67 12126 -67 4 xa[6]
port 138 nsew
rlabel metal2 s 12391 -67 12391 -67 4 xa[5]
port 139 nsew
rlabel metal2 s 12656 -67 12656 -67 4 xa[4]
port 140 nsew
rlabel metal2 s 13713 -67 13713 -67 4 xa[0]
port 141 nsew
rlabel metal2 s 6038 31 6038 31 4 men
port 142 nsew
rlabel metal2 s 12919 -67 12919 -67 4 xa[3]
port 143 nsew
rlabel metal2 s 13184 -67 13184 -67 4 xa[2]
port 144 nsew
rlabel metal2 s 13449 -67 13449 -67 4 xa[1]
port 145 nsew
rlabel metal2 s 9298 -67 9298 -67 4 xc[0]
port 146 nsew
rlabel metal2 s 9034 -67 9034 -67 4 xc[1]
port 147 nsew
rlabel metal3 s 44 927 44 927 4 LWL[1]
port 91 nsew
rlabel metal3 s 44 310 44 310 4 LWL[0]
port 92 nsew
rlabel metal3 s 44 1522 44 1522 4 LWL[2]
port 90 nsew
rlabel metal3 s 44 2138 44 2138 4 LWL[3]
port 89 nsew
rlabel metal3 s 44 2732 44 2732 4 LWL[4]
port 88 nsew
rlabel metal3 s 44 3348 44 3348 4 LWL[5]
port 87 nsew
rlabel metal3 s 44 3946 44 3946 4 LWL[6]
port 95 nsew
rlabel metal3 s 44 4562 44 4562 4 LWL[7]
port 97 nsew
rlabel metal3 s 44 5158 44 5158 4 LWL[8]
port 93 nsew
rlabel metal3 s 44 5774 44 5774 4 LWL[9]
port 94 nsew
rlabel metal3 s 44 6370 44 6370 4 LWL[10]
port 78 nsew
rlabel metal3 s 44 6986 44 6986 4 LWL[11]
port 79 nsew
rlabel metal3 s 44 7581 44 7581 4 LWL[12]
port 80 nsew
rlabel metal3 s 44 8197 44 8197 4 LWL[13]
port 81 nsew
rlabel metal3 s 44 8794 44 8794 4 LWL[14]
port 82 nsew
rlabel metal3 s 44 9410 44 9410 4 LWL[15]
port 83 nsew
rlabel metal3 s 44 10006 44 10006 4 LWL[16]
port 84 nsew
rlabel metal3 s 44 10622 44 10622 4 LWL[17]
port 85 nsew
rlabel metal3 s 44 11218 44 11218 4 LWL[18]
port 86 nsew
rlabel metal3 s 44 11834 44 11834 4 LWL[19]
port 68 nsew
rlabel metal3 s 44 13046 44 13046 4 LWL[21]
port 70 nsew
rlabel metal3 s 44 12430 44 12430 4 LWL[20]
port 69 nsew
rlabel metal3 s 44 13642 44 13642 4 LWL[22]
port 71 nsew
rlabel metal3 s 44 14258 44 14258 4 LWL[23]
port 72 nsew
rlabel metal3 s 44 14854 44 14854 4 LWL[24]
port 73 nsew
rlabel metal3 s 44 15470 44 15470 4 LWL[25]
port 74 nsew
rlabel metal3 s 44 16062 44 16062 4 LWL[26]
port 75 nsew
rlabel metal3 s 44 16678 44 16678 4 LWL[27]
port 76 nsew
rlabel metal3 s 44 18488 44 18488 4 LWL[30]
port 99 nsew
rlabel metal3 s 44 17894 44 17894 4 LWL[29]
port 98 nsew
rlabel metal3 s 44 17278 44 17278 4 LWL[28]
port 77 nsew
rlabel metal3 s 44 19106 44 19106 4 LWL[31]
port 67 nsew
rlabel metal3 s 44 21531 44 21531 4 LWL[35]
port 61 nsew
rlabel metal3 s 44 20912 44 20912 4 LWL[34]
port 62 nsew
rlabel metal3 s 44 20320 44 20320 4 LWL[33]
port 63 nsew
rlabel metal3 s 44 19700 44 19700 4 LWL[32]
port 96 nsew
rlabel metal3 s 44 22124 44 22124 4 LWL[36]
port 60 nsew
rlabel metal3 s 44 22743 44 22743 4 LWL[37]
port 59 nsew
rlabel metal3 s 44 23336 44 23336 4 LWL[38]
port 58 nsew
rlabel metal3 s 44 23955 44 23955 4 LWL[39]
port 57 nsew
rlabel metal3 s 44 24549 44 24549 4 LWL[40]
port 56 nsew
rlabel metal3 s 44 25166 44 25166 4 LWL[41]
port 55 nsew
rlabel metal3 s 44 25761 44 25761 4 LWL[42]
port 54 nsew
rlabel metal3 s 44 26380 44 26380 4 LWL[43]
port 53 nsew
rlabel metal3 s 44 26973 44 26973 4 LWL[44]
port 52 nsew
rlabel metal3 s 44 27591 44 27591 4 LWL[45]
port 51 nsew
rlabel metal3 s 44 28185 44 28185 4 LWL[46]
port 50 nsew
rlabel metal3 s 44 28803 44 28803 4 LWL[47]
port 49 nsew
rlabel metal3 s 44 29397 44 29397 4 LWL[48]
port 48 nsew
rlabel metal3 s 44 30016 44 30016 4 LWL[49]
port 47 nsew
rlabel metal3 s 44 30609 44 30609 4 LWL[50]
port 46 nsew
rlabel metal3 s 44 31228 44 31228 4 LWL[51]
port 45 nsew
rlabel metal3 s 44 31821 44 31821 4 LWL[52]
port 44 nsew
rlabel metal3 s 44 32440 44 32440 4 LWL[53]
port 43 nsew
rlabel metal3 s 44 33033 44 33033 4 LWL[54]
port 42 nsew
rlabel metal3 s 44 33651 44 33651 4 LWL[55]
port 41 nsew
rlabel metal3 s 44 34245 44 34245 4 LWL[56]
port 40 nsew
rlabel metal3 s 44 34863 44 34863 4 LWL[57]
port 39 nsew
rlabel metal3 s 44 35457 44 35457 4 LWL[58]
port 38 nsew
rlabel metal3 s 44 36075 44 36075 4 LWL[59]
port 37 nsew
rlabel metal3 s 44 36668 44 36668 4 LWL[60]
port 36 nsew
rlabel metal3 s 44 37497 44 37497 4 LWL[61]
port 35 nsew
rlabel metal3 s 44 38091 44 38091 4 LWL[62]
port 34 nsew
rlabel metal3 s 93 38801 93 38801 4 vdd
port 65 nsew
rlabel metal3 s 35 38506 35 38506 4 LWL[63]
port 33 nsew
rlabel metal3 s 472 39092 472 39092 4 DLWL
port 66 nsew
rlabel metal3 s 19393 928 19393 928 4 RWL[1]
port 116 nsew
rlabel metal3 s 19393 312 19393 312 4 RWL[0]
port 115 nsew
rlabel metal3 s 19393 1522 19393 1522 4 RWL[2]
port 114 nsew
rlabel metal3 s 19393 2138 19393 2138 4 RWL[3]
port 117 nsew
rlabel metal3 s 19393 2732 19393 2732 4 RWL[4]
port 113 nsew
rlabel metal3 s 19393 3348 19393 3348 4 RWL[5]
port 118 nsew
rlabel metal3 s 19393 3946 19393 3946 4 RWL[6]
port 112 nsew
rlabel metal3 s 19393 4562 19393 4562 4 RWL[7]
port 119 nsew
rlabel metal3 s 19393 5158 19393 5158 4 RWL[8]
port 120 nsew
rlabel metal3 s 19393 5774 19393 5774 4 RWL[9]
port 121 nsew
rlabel metal3 s 19393 6370 19393 6370 4 RWL[10]
port 122 nsew
rlabel metal3 s 19393 6986 19393 6986 4 RWL[11]
port 123 nsew
rlabel metal3 s 19393 7582 19393 7582 4 RWL[12]
port 124 nsew
rlabel metal3 s 19393 8198 19393 8198 4 RWL[13]
port 125 nsew
rlabel metal3 s 19393 8794 19393 8794 4 RWL[14]
port 126 nsew
rlabel metal3 s 19393 9410 19393 9410 4 RWL[15]
port 127 nsew
rlabel metal3 s 19393 10006 19393 10006 4 RWL[16]
port 128 nsew
rlabel metal3 s 19393 10622 19393 10622 4 RWL[17]
port 129 nsew
rlabel metal3 s 19393 11218 19393 11218 4 RWL[18]
port 130 nsew
rlabel metal3 s 19393 11834 19393 11834 4 RWL[19]
port 131 nsew
rlabel metal3 s 19393 13046 19393 13046 4 RWL[21]
port 111 nsew
rlabel metal3 s 19393 12430 19393 12430 4 RWL[20]
port 132 nsew
rlabel metal3 s 19393 13642 19393 13642 4 RWL[22]
port 110 nsew
rlabel metal3 s 19393 14258 19393 14258 4 RWL[23]
port 109 nsew
rlabel metal3 s 19393 15470 19393 15470 4 RWL[25]
port 107 nsew
rlabel metal3 s 19393 14854 19393 14854 4 RWL[24]
port 108 nsew
rlabel metal3 s 19393 16682 19393 16682 4 RWL[27]
port 105 nsew
rlabel metal3 s 19393 16066 19393 16066 4 RWL[26]
port 106 nsew
rlabel metal3 s 19393 17894 19393 17894 4 RWL[29]
port 103 nsew
rlabel metal3 s 19393 17278 19393 17278 4 RWL[28]
port 104 nsew
rlabel metal3 s 19393 19106 19393 19106 4 RWL[31]
port 101 nsew
rlabel metal3 s 19393 18490 19393 18490 4 RWL[30]
port 102 nsew
rlabel metal3 s 19393 19699 19393 19699 4 RWL[32]
port 100 nsew
rlabel metal3 s 19393 20319 19393 20319 4 RWL[33]
port 2 nsew
rlabel metal3 s 19393 20913 19393 20913 4 RWL[34]
port 3 nsew
rlabel metal3 s 19393 21531 19393 21531 4 RWL[35]
port 4 nsew
rlabel metal3 s 19393 22124 19393 22124 4 RWL[36]
port 5 nsew
rlabel metal3 s 19393 22743 19393 22743 4 RWL[37]
port 6 nsew
rlabel metal3 s 19393 23337 19393 23337 4 RWL[38]
port 7 nsew
rlabel metal3 s 19393 23955 19393 23955 4 RWL[39]
port 8 nsew
rlabel metal3 s 19393 24549 19393 24549 4 RWL[40]
port 9 nsew
rlabel metal3 s 19393 25167 19393 25167 4 RWL[41]
port 10 nsew
rlabel metal3 s 19393 25761 19393 25761 4 RWL[42]
port 11 nsew
rlabel metal3 s 19393 26379 19393 26379 4 RWL[43]
port 12 nsew
rlabel metal3 s 19393 26973 19393 26973 4 RWL[44]
port 13 nsew
rlabel metal3 s 19393 27592 19393 27592 4 RWL[45]
port 14 nsew
rlabel metal3 s 19393 28186 19393 28186 4 RWL[46]
port 15 nsew
rlabel metal3 s 19393 28803 19393 28803 4 RWL[47]
port 16 nsew
rlabel metal3 s 19392 29398 19392 29398 4 RWL[48]
port 17 nsew
rlabel metal3 s 19392 30016 19392 30016 4 RWL[49]
port 18 nsew
rlabel metal3 s 19392 30609 19392 30609 4 RWL[50]
port 19 nsew
rlabel metal3 s 19392 31227 19392 31227 4 RWL[51]
port 20 nsew
rlabel metal3 s 19392 31821 19392 31821 4 RWL[52]
port 21 nsew
rlabel metal3 s 19392 32439 19392 32439 4 RWL[53]
port 22 nsew
rlabel metal3 s 19392 33033 19392 33033 4 RWL[54]
port 23 nsew
rlabel metal3 s 19392 33651 19392 33651 4 RWL[55]
port 24 nsew
rlabel metal3 s 19392 34245 19392 34245 4 RWL[56]
port 25 nsew
rlabel metal3 s 19392 34863 19392 34863 4 RWL[57]
port 26 nsew
rlabel metal3 s 19392 35457 19392 35457 4 RWL[58]
port 27 nsew
rlabel metal3 s 19392 36075 19392 36075 4 RWL[59]
port 28 nsew
rlabel metal3 s 19392 36669 19392 36669 4 RWL[60]
port 29 nsew
rlabel metal3 s 19392 37287 19392 37287 4 RWL[61]
port 30 nsew
rlabel metal3 s 19392 37881 19392 37881 4 RWL[62]
port 31 nsew
rlabel metal3 s 19392 38499 19392 38499 4 RWL[63]
port 32 nsew
rlabel metal3 s 18968 39092 18968 39092 4 DRWL
port 1 nsew
rlabel metal3 s 93 39401 93 39401 4 vss
port 64 nsew
<< end >>
