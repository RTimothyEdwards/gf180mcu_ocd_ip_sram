magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal2 >>
rect -118 101 119 118
rect -118 -181 -102 101
rect 102 -181 119 101
rect -118 -198 119 -181
<< via2 >>
rect -102 -181 102 101
<< metal3 >>
rect -119 101 119 118
rect -119 -181 -102 101
rect 102 -181 119 101
rect -119 -198 119 -181
<< end >>
