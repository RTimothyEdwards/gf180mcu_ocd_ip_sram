magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nmos >>
rect 0 0 56 614
<< ndiff >>
rect -88 601 0 614
rect -88 13 -75 601
rect -29 13 0 601
rect -88 0 0 13
rect 56 601 144 614
rect 56 13 85 601
rect 131 13 144 601
rect 56 0 144 13
<< ndiffc >>
rect -75 13 -29 601
rect 85 13 131 601
<< polysilicon >>
rect 0 614 56 658
rect 0 -44 56 0
<< metal1 >>
rect -75 601 -29 614
rect -75 0 -29 13
rect 85 601 131 614
rect 85 0 131 13
<< labels >>
flabel ndiffc -40 307 -40 307 0 FreeSans 93 0 0 0 S
flabel ndiffc 96 307 96 307 0 FreeSans 93 0 0 0 D
<< end >>
