magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal2 >>
rect -119 713 119 732
rect -119 -713 -102 713
rect 102 -713 119 713
rect -119 -732 119 -713
<< via2 >>
rect -102 -713 102 713
<< metal3 >>
rect -119 713 119 732
rect -119 -713 -102 713
rect 102 -713 119 713
rect -119 -732 119 -713
<< end >>
