magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -44 409 44 427
rect -44 -409 -28 409
rect 28 -409 44 409
rect -44 -427 44 -409
<< via2 >>
rect -28 -409 28 409
<< metal3 >>
rect -45 409 45 427
rect -45 -409 -28 409
rect 28 -409 45 409
rect -45 -427 45 -409
<< end >>
