magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< nwell >>
rect 1546 3720 3253 4738
rect 1521 3402 3287 3720
rect 1970 901 3163 974
<< psubdiff >>
rect 1395 4897 3523 5013
rect 3412 1216 3523 4897
rect 3412 762 3445 1216
rect 3491 762 3523 1216
rect 1727 694 1838 734
rect 1727 693 1839 694
rect 3412 693 3523 762
rect 1727 578 3523 693
<< psubdiffcont >>
rect 3445 762 3491 1216
<< polysilicon >>
rect 2217 4691 2594 4761
rect 2217 4576 2273 4691
rect 2377 4576 2433 4691
rect 2538 4576 2594 4691
rect 1734 4076 1790 4291
rect 1894 4076 1950 4291
rect 2380 4076 2436 4291
rect 2844 4076 2900 4291
rect 3004 4076 3060 4291
rect 1466 3745 1951 3784
rect 2844 3745 3303 3784
rect 1939 3399 2003 3458
rect 1784 3242 1873 3308
rect 1784 2934 1841 3242
rect 2107 3161 2164 3459
rect 2107 3126 2186 3161
rect 1944 3090 2186 3126
rect 1944 3080 2162 3090
rect 1944 2934 2000 3080
rect 2105 2934 2162 3080
rect 2271 2994 2324 3467
rect 2440 3465 2486 3467
rect 2266 2934 2324 2994
rect 2428 3316 2486 3465
rect 2428 3245 2530 3316
rect 2428 2934 2484 3245
rect 2588 3126 2646 3467
rect 2750 3407 2884 3466
rect 2886 3238 2967 3308
rect 2588 3078 2806 3126
rect 2588 2934 2644 3078
rect 2749 2995 2806 3078
rect 2750 2934 2806 2995
rect 2909 2934 2967 3238
rect 3071 2444 3127 2547
rect 1813 2042 1869 2046
rect 1973 2042 2029 2046
rect 2135 2042 2191 2046
rect 2295 2042 2351 2046
rect 2457 2042 2513 2046
rect 2617 2042 2673 2046
rect 2779 2042 2835 2046
rect 2939 2042 2995 2046
rect 1812 2034 2995 2042
rect 1812 1946 2993 2034
rect 2139 1451 2195 1589
rect 2120 1379 2355 1451
rect 2139 1302 2195 1379
rect 2299 1302 2355 1379
rect 2460 1302 2516 1589
rect 2620 1568 2677 1589
rect 2781 1568 2837 1589
rect 2620 1527 2837 1568
rect 2620 1451 2676 1527
rect 2590 1379 2676 1451
rect 2941 1415 2997 1589
rect 2620 1302 2676 1379
rect 2781 1370 2997 1415
rect 2781 1302 2837 1370
rect 2941 1302 2997 1370
<< metal1 >>
rect 1229 5555 1817 5623
rect 1752 5476 1817 5555
rect 2153 5545 3150 5613
rect 1752 5408 3150 5476
rect 1229 5234 3419 5331
rect 875 5085 3150 5153
rect 1291 4904 3517 5007
rect 2289 4803 2526 4856
rect 1290 1895 1390 4748
rect 1670 4696 2317 4748
rect 1670 4322 1720 4696
rect 1979 4323 2025 4696
rect 2267 4328 2317 4696
rect 2371 4689 2437 4803
rect 2491 4696 3138 4748
rect 2491 4328 2541 4696
rect 2757 4328 2838 4696
rect 3087 4328 3138 4696
rect 1985 4322 2018 4323
rect 1664 4148 1726 4272
rect 1990 4148 2053 4272
rect 2294 4207 3141 4272
rect 1664 4089 2513 4148
rect 1663 4083 2513 4089
rect 1663 3852 1726 4083
rect 1444 2036 1495 3798
rect 1819 3776 1865 3887
rect 1985 3826 2033 4083
rect 2302 3776 2354 3909
rect 2767 3900 2814 4207
rect 1713 3724 2354 3776
rect 2465 3776 2517 3900
rect 2781 3899 2814 3900
rect 2927 3776 2979 3892
rect 3089 3853 3141 4207
rect 3095 3852 3127 3853
rect 2465 3724 3038 3776
rect 3250 3751 3441 3798
rect 1600 3656 1666 3657
rect 1584 3443 1666 3656
rect 1632 3041 1682 3163
rect 1713 3098 1764 3724
rect 2205 3656 2271 3657
rect 2536 3656 2601 3657
rect 1875 3404 1955 3622
rect 1632 2989 1757 3041
rect 1707 2893 1757 2989
rect 2029 2896 2082 3626
rect 2200 3443 2282 3656
rect 2158 3236 2327 3320
rect 2158 3081 2305 3168
rect 2375 3043 2425 3622
rect 2527 3443 2607 3656
rect 2477 3236 2630 3320
rect 2503 3081 2657 3168
rect 2350 2990 2425 3043
rect 2720 3038 2770 3621
rect 2827 3404 2908 3628
rect 2886 3245 2940 3312
rect 2987 3098 3038 3724
rect 3092 3656 3158 3657
rect 3092 3443 3173 3656
rect 3132 3165 3182 3313
rect 3131 3097 3182 3165
rect 3132 3041 3182 3097
rect 2350 2893 2400 2990
rect 2674 2984 2770 3038
rect 2996 2989 3182 3041
rect 2674 2893 2720 2984
rect 2996 2893 3042 2989
rect 1549 2447 1630 2893
rect 1875 2531 1955 2647
rect 2200 2531 2282 2647
rect 2527 2531 2607 2647
rect 2834 2531 2881 2647
rect 1875 2466 2881 2531
rect 1892 2092 1972 2466
rect 2205 2092 2286 2466
rect 2519 2092 2599 2466
rect 2832 2092 2913 2466
rect 3178 2447 3259 2896
rect 3390 2036 3441 3751
rect 1444 1952 3441 2036
rect 1290 1795 1831 1895
rect 1290 1792 1833 1795
rect 1733 687 1833 1792
rect 2224 1439 2270 1637
rect 2224 1391 2590 1439
rect 2047 859 2128 1261
rect 2224 1235 2270 1391
rect 2361 859 2441 1261
rect 2674 859 2755 1261
rect 2987 859 3068 1261
rect 3418 1216 3517 1278
rect 3418 762 3445 1216
rect 3491 762 3517 1216
rect 3418 687 3517 762
rect 1733 584 3517 687
<< metal2 >>
rect 1754 5623 1816 5702
rect 2146 5623 2208 5734
rect 1702 5613 1816 5623
rect 1702 5555 1765 5613
rect 2135 5555 2208 5623
rect 1968 5408 2034 5476
rect 2659 5408 2722 5702
rect 3053 5613 3116 5747
rect 2795 5545 3116 5613
rect 1969 4748 2034 5408
rect 1968 4696 2034 4748
rect 2371 4689 2437 5153
rect 2795 4680 2860 5545
rect 1816 4272 1879 4554
rect 1449 4207 1879 4272
rect 1449 3313 1512 4207
rect 2293 4083 2359 4350
rect 2451 4083 2517 4350
rect 2926 4274 2991 4554
rect 2926 4206 3287 4274
rect 1449 3245 3122 3313
rect 1449 1946 1512 3245
rect 3221 3165 3287 4206
rect 1671 3097 3287 3165
rect 3221 1947 3287 3097
rect 1449 1881 1986 1946
rect 1924 1382 1986 1881
rect 2995 1879 3434 1947
rect 2370 1576 2435 1751
rect 2678 1576 2744 1751
rect 2992 1576 3058 1751
rect 2370 1508 2744 1576
rect 2842 1508 3058 1576
rect 2520 376 2586 1508
rect 2842 393 2907 1508
rect 3126 1382 3192 1879
<< metal3 >>
rect 1701 5545 2191 5613
rect 1701 5476 1766 5545
rect 1178 5408 1766 5476
rect -249 3068 3468 4974
rect -249 1011 3504 2867
rect -249 385 3504 886
use M1_NWELL06_256x8m81  M1_NWELL06_256x8m81_0
timestamp 1763564386
transform 1 0 2566 0 1 900
box -596 -159 597 159
use M1_NWELL_01_R90_256x8m81  M1_NWELL_01_R90_256x8m81_0
timestamp 1763564386
transform 0 -1 1619 1 0 3561
box -159 -154 159 154
use M1_NWELL_01_R90_256x8m81  M1_NWELL_01_R90_256x8m81_1
timestamp 1763564386
transform 0 -1 3132 1 0 3561
box -159 -154 159 154
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_0
timestamp 1763564386
transform -1 0 2720 0 1 1994
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_1
timestamp 1763564386
transform -1 0 2925 0 1 1994
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_2
timestamp 1763564386
transform 1 0 3154 0 1 2492
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_3
timestamp 1763564386
transform -1 0 2092 0 1 1994
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_4
timestamp 1763564386
transform 1 0 1647 0 1 2491
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_5
timestamp 1763564386
transform 1 0 1880 0 1 1994
box -67 -48 67 47
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_6
timestamp 1763564386
transform -1 0 2404 0 1 1994
box -67 -48 67 47
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_0
timestamp 1763564386
transform 1 0 2296 0 1 3278
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_1
timestamp 1763564386
transform 1 0 2181 0 1 3127
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_2
timestamp 1763564386
transform 1 0 1918 0 1 3428
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_3
timestamp 1763564386
transform 1 0 1495 0 1 3775
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_4
timestamp 1763564386
transform 1 0 1902 0 1 3278
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_5
timestamp 1763564386
transform 1 0 2633 0 1 3127
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_6
timestamp 1763564386
transform 1 0 2501 0 1 3278
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_7
timestamp 1763564386
transform 1 0 2906 0 1 3278
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_8
timestamp 1763564386
transform 1 0 2855 0 1 3430
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_9
timestamp 1763564386
transform 1 0 3273 0 1 3775
box -36 -36 36 36
use M1_POLY24310591302031_256x8m81  M1_POLY24310591302031_256x8m81_10
timestamp 1763564386
transform 1 0 2404 0 1 4731
box -36 -36 36 36
use M1_POLY24310591302033_256x8m81  M1_POLY24310591302033_256x8m81_0
timestamp 1763564386
transform 1 0 2533 0 1 1415
box -62 -36 62 36
use M1_POLY24310591302033_256x8m81  M1_POLY24310591302033_256x8m81_1
timestamp 1763564386
transform 1 0 3052 0 1 1407
box -62 -36 62 36
use M1_POLY24310591302033_256x8m81  M1_POLY24310591302033_256x8m81_2
timestamp 1763564386
transform 1 0 2071 0 1 1415
box -62 -36 62 36
use M1_PSUB$$46555180_256x8m81  M1_PSUB$$46555180_256x8m81_0
timestamp 1763564386
transform 1 0 2407 0 1 4956
box -996 -58 996 57
use M1_PSUB$$46556204_256x8m81  M1_PSUB$$46556204_256x8m81_0
timestamp 1763564386
transform 1 0 1340 0 1 3515
box -56 -1729 56 1498
use M1_PSUB$$46557228_256x8m81  M1_PSUB$$46557228_256x8m81_0
timestamp 1763564386
transform 1 0 1561 0 1 1844
box -277 -58 277 58
use M1_PSUB$$46558252_256x8m81  M1_PSUB$$46558252_256x8m81_0
timestamp 1763564386
transform 1 0 2571 0 1 636
box -665 -58 665 57
use M1_PSUB_04_R90_256x8m81  M1_PSUB_04_R90_256x8m81_0
timestamp 1763564386
transform 0 -1 1782 1 0 1051
box -461 -56 571 55
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_0
timestamp 1763564386
transform 1 0 3035 0 1 2484
box -119 -46 119 46
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_1
timestamp 1763564386
transform 1 0 1769 0 1 2484
box -119 -46 119 46
use nmos_1p2$$45107244_256x8m81  nmos_1p2$$45107244_256x8m81_0
timestamp 1763564386
transform -1 0 2900 0 -1 1839
box -185 -44 527 255
use nmos_1p2$$46550060_256x8m81  nmos_1p2$$46550060_256x8m81_0
timestamp 1763564386
transform 1 0 2024 0 1 2087
box -299 -44 1060 309
use nmos_1p2$$46551084_256x8m81  nmos_1p2$$46551084_256x8m81_0
timestamp 1763564386
transform -1 0 2181 0 -1 1839
box -102 -44 130 255
use nmos_1p2$$46552108_256x8m81  nmos_1p2$$46552108_256x8m81_0
timestamp 1763564386
transform 1 0 1996 0 1 2581
box -301 -45 1060 363
use nmos_1p2$$46553132_256x8m81  nmos_1p2$$46553132_256x8m81_0
timestamp 1763564386
transform 1 0 3085 0 1 2581
box -102 -44 130 362
use nmos_1p2$$46553132_256x8m81  nmos_1p2$$46553132_256x8m81_1
timestamp 1763564386
transform 1 0 1638 0 1 2581
box -102 -44 130 362
use pmos_1p2$$46285868_256x8m81  pmos_1p2$$46285868_256x8m81_0
timestamp 1763564386
transform 1 0 2394 0 1 3826
box -188 -86 216 297
use pmos_1p2$$46286892_256x8m81  pmos_1p2$$46286892_256x8m81_0
timestamp 1763564386
transform 1 0 2287 0 1 4322
box -244 -86 481 297
use pmos_1p2$$46549036_256x8m81  pmos_1p2$$46549036_256x8m81_0
timestamp 1763564386
transform -1 0 2843 0 -1 1261
box -328 -86 878 297
use pmos_1p2$$46896172_256x8m81  pmos_1p2$$46896172_256x8m81_0
timestamp 1763564386
transform 1 0 2206 0 1 3501
box -272 -86 613 170
use pmos_1p2$$46897196_256x8m81  pmos_1p2$$46897196_256x8m81_0
timestamp 1763564386
transform 1 0 1776 0 1 4322
box -216 -86 348 297
use pmos_1p2$$46897196_256x8m81  pmos_1p2$$46897196_256x8m81_1
timestamp 1763564386
transform 1 0 1776 0 1 3826
box -216 -86 348 297
use pmos_1p2$$46897196_256x8m81  pmos_1p2$$46897196_256x8m81_2
timestamp 1763564386
transform 1 0 2886 0 1 4322
box -216 -86 348 297
use pmos_1p2$$46897196_256x8m81  pmos_1p2$$46897196_256x8m81_3
timestamp 1763564386
transform 1 0 2886 0 1 3826
box -216 -86 348 297
use pmos_1p2$$46898220_256x8m81  pmos_1p2$$46898220_256x8m81_0
timestamp 1763564386
transform 1 0 1962 0 1 3501
box -188 -86 216 170
use pmos_1p2$$46898220_256x8m81  pmos_1p2$$46898220_256x8m81_1
timestamp 1763564386
transform 1 0 2763 0 1 3501
box -188 -86 216 170
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_0
timestamp 1763564386
transform 1 0 3436 0 1 1058
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_1
timestamp 1763564386
transform 1 0 2683 0 1 2164
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_2
timestamp 1763564386
transform -1 0 2590 0 -1 1870
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_3
timestamp 1763564386
transform -1 0 2902 0 -1 1870
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_4
timestamp 1763564386
transform 1 0 2989 0 1 2164
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_5
timestamp 1763564386
transform 1 0 2370 0 1 2164
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_6
timestamp 1763564386
transform -1 0 2123 0 -1 1750
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_7
timestamp 1763564386
transform 1 0 1766 0 1 1058
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_8
timestamp 1763564386
transform 1 0 1766 0 1 1471
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_9
timestamp 1763564386
transform 1 0 1750 0 1 2164
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_10
timestamp 1763564386
transform 1 0 2056 0 1 2164
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_11
timestamp 1763564386
transform 1 0 1890 0 1 3405
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_12
timestamp 1763564386
transform 1 0 2205 0 1 3445
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_13
timestamp 1763564386
transform 1 0 1592 0 1 3445
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_14
timestamp 1763564386
transform 1 0 2135 0 1 4387
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_15
timestamp 1763564386
transform 1 0 2536 0 1 3445
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_16
timestamp 1763564386
transform 1 0 2605 0 1 4387
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_17
timestamp 1763564386
transform 1 0 2828 0 1 3405
box -9 0 73 215
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_18
timestamp 1763564386
transform 1 0 3092 0 1 3445
box -9 0 73 215
use via1_2_x2_R90_256x8m81  via1_2_x2_R90_256x8m81_0
timestamp 1763564386
transform 0 -1 2281 1 0 5545
box -9 0 73 215
use via1_2_x2_R270_256x8m81  via1_2_x2_R270_256x8m81_0
timestamp 1763564386
transform 0 1 2983 -1 0 910
box -9 0 75 215
use via1_2_x2_R270_256x8m81  via1_2_x2_R270_256x8m81_1
timestamp 1763564386
transform 0 1 1906 -1 0 910
box -9 0 75 215
use via1_2_x2_R270_256x8m81  via1_2_x2_R270_256x8m81_2
timestamp 1763564386
transform 0 1 2227 -1 0 910
box -9 0 75 215
use via1_256x8m81  via1_256x8m81_0
timestamp 1763564386
transform 1 0 2371 0 -1 4783
box 0 0 65 92
use via1_R90_256x8m81  via1_R90_256x8m81_0
timestamp 1763564386
transform 0 -1 3154 1 0 2464
box 0 0 65 89
use via1_R90_256x8m81  via1_R90_256x8m81_1
timestamp 1763564386
transform 0 -1 1740 1 0 2464
box 0 0 65 89
use via1_R90_256x8m81  via1_R90_256x8m81_2
timestamp 1763564386
transform 0 -1 1764 1 0 3098
box 0 0 65 89
use via1_R90_256x8m81  via1_R90_256x8m81_3
timestamp 1763564386
transform 0 -1 3077 1 0 3245
box 0 0 65 89
use via1_R90_256x8m81  via1_R90_256x8m81_4
timestamp 1763564386
transform 0 -1 3197 1 0 3098
box 0 0 65 89
use via1_R90_256x8m81  via1_R90_256x8m81_5
timestamp 1763564386
transform 0 -1 2516 1 0 4084
box 0 0 65 89
use via1_R90_256x8m81  via1_R90_256x8m81_6
timestamp 1763564386
transform 0 1 2293 1 0 4204
box 0 0 65 89
use via1_R270_256x8m81  via1_R270_256x8m81_0
timestamp 1763564386
transform 0 -1 2047 -1 0 4763
box 0 0 67 89
use via1_R270_256x8m81  via1_R270_256x8m81_1
timestamp 1763564386
transform 0 1 2158 -1 0 3164
box 0 0 67 89
use via1_R270_256x8m81  via1_R270_256x8m81_2
timestamp 1763564386
transform 0 1 2235 -1 0 3312
box 0 0 67 89
use via1_R270_256x8m81  via1_R270_256x8m81_3
timestamp 1763564386
transform 0 -1 2450 -1 0 5152
box 0 0 67 89
use via1_R270_256x8m81  via1_R270_256x8m81_4
timestamp 1763564386
transform 0 -1 2842 -1 0 4748
box 0 0 67 89
use via1_R270_256x8m81  via1_R270_256x8m81_5
timestamp 1763564386
transform 0 1 2561 -1 0 3164
box 0 0 67 89
use via1_R270_256x8m81  via1_R270_256x8m81_6
timestamp 1763564386
transform 0 1 2359 -1 0 3164
box 0 0 67 89
use via1_R270_256x8m81  via1_R270_256x8m81_7
timestamp 1763564386
transform 0 1 2484 -1 0 3312
box 0 0 67 89
use via1_x2_256x8m81  via1_x2_256x8m81_0
timestamp 1763564386
transform -1 0 2907 0 1 1042
box -8 0 72 222
use via1_x2_256x8m81  via1_x2_256x8m81_1
timestamp 1763564386
transform 1 0 2993 0 1 1528
box -8 0 72 222
use via1_x2_256x8m81  via1_x2_256x8m81_2
timestamp 1763564386
transform 1 0 2520 0 1 1042
box -8 0 72 222
use via1_x2_256x8m81  via1_x2_256x8m81_3
timestamp 1763564386
transform -1 0 2744 0 1 1528
box -8 0 72 222
use via1_x2_256x8m81  via1_x2_256x8m81_4
timestamp 1763564386
transform -1 0 2434 0 1 1528
box -8 0 72 222
use via1_x2_256x8m81  via1_x2_256x8m81_5
timestamp 1763564386
transform 1 0 1817 0 1 4332
box -8 0 72 222
use via1_x2_256x8m81  via1_x2_256x8m81_6
timestamp 1763564386
transform 1 0 2926 0 1 4332
box -8 0 72 222
use via1_x2_256x8m81  via1_x2_256x8m81_7
timestamp 1763564386
transform 1 0 2452 0 1 4332
box -8 0 72 222
use via1_x2_256x8m81  via1_x2_256x8m81_8
timestamp 1763564386
transform -1 0 2358 0 1 4332
box -8 0 72 222
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_0
timestamp 1763564386
transform 0 -1 3191 1 0 1375
box -8 0 72 215
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_1
timestamp 1763564386
transform 0 -1 2139 1 0 1383
box -8 0 72 215
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_2
timestamp 1763564386
transform 0 -1 2110 1 0 5407
box -8 0 72 215
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_3
timestamp 1763564386
transform 0 -1 1843 1 0 5555
box -8 0 72 215
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_4
timestamp 1763564386
transform 0 -1 2713 1 0 5409
box -8 0 72 215
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_5
timestamp 1763564386
transform 0 -1 3147 1 0 5545
box -8 0 72 215
use via1_x2_R270_256x8m81  via1_x2_R270_256x8m81_0
timestamp 1763564386
transform 0 1 1878 -1 0 3312
box -8 0 75 215
use via1_x2_R270_256x8m81  via1_x2_R270_256x8m81_1
timestamp 1763564386
transform 0 1 2718 -1 0 3312
box -8 0 75 215
use via2_x2_R90_256x8m81  via2_x2_R90_256x8m81_0
timestamp 1763564386
transform 0 -1 1394 1 0 5409
box -9 0 73 215
<< labels >>
rlabel metal2 s 2007 4921 2007 4921 4 d
port 5 nsew
rlabel metal1 s 2416 5285 2416 5285 4 wep
port 7 nsew
rlabel metal1 s 1428 5106 1428 5106 4 pcb
port 9 nsew
rlabel metal1 s 2402 5446 2402 5446 4 d
port 5 nsew
rlabel metal2 s 2826 4921 2826 4921 4 db
port 4 nsew
rlabel metal1 s 2405 5587 2405 5587 4 db
port 4 nsew
rlabel metal3 s 722 646 722 646 4 vdd
port 1 nsew
rlabel metal1 s 3129 2012 3129 2012 4 se
port 8 nsew
rlabel metal3 s 872 2017 872 2017 4 vss
port 2 nsew
rlabel metal2 s 2877 435 2877 435 4 qn
port 6 nsew
rlabel metal2 s 2553 435 2553 435 4 qp
port 3 nsew
<< end >>
