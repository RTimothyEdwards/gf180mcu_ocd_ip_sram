magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< metal2 >>
rect -99 92 99 99
rect -99 -92 -92 92
rect 92 -92 99 92
rect -99 -99 99 -92
<< via2 >>
rect -92 -92 92 92
<< metal3 >>
rect -99 92 99 99
rect -99 -92 -92 92
rect 92 -92 99 92
rect -99 -99 99 -92
<< end >>
