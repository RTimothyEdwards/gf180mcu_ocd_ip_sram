magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -44 257 44 275
rect -44 -87 -28 257
rect 28 -87 44 257
rect -44 -105 44 -87
<< via2 >>
rect -28 -87 28 257
<< metal3 >>
rect -45 257 45 275
rect -45 -87 -28 257
rect 28 -87 45 257
rect -45 -105 45 -87
<< end >>
