magic
tech gf180mcuD
magscale 1 10
timestamp 1765482800
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_0
timestamp 1764626446
transform -1 0 668 0 1 18896
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_1
timestamp 1764626446
transform -1 0 668 0 1 38288
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_2
timestamp 1764626446
transform -1 0 668 0 1 716
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_3
timestamp 1764626446
transform -1 0 668 0 1 3140
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_4
timestamp 1764626446
transform -1 0 668 0 1 4352
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_5
timestamp 1764626446
transform -1 0 668 0 1 5564
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_6
timestamp 1764626446
transform -1 0 668 0 1 6776
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_7
timestamp 1764626446
transform -1 0 668 0 1 7988
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_8
timestamp 1764626446
transform -1 0 668 0 1 9200
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_9
timestamp 1764626446
transform -1 0 668 0 1 10412
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_10
timestamp 1764626446
transform -1 0 668 0 1 11624
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_11
timestamp 1764626446
transform -1 0 668 0 1 12836
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_12
timestamp 1764626446
transform -1 0 668 0 1 14048
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_13
timestamp 1764626446
transform -1 0 668 0 1 15260
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_14
timestamp 1764626446
transform -1 0 668 0 1 16472
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_15
timestamp 1764626446
transform -1 0 668 0 1 17684
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_16
timestamp 1764626446
transform -1 0 668 0 1 21320
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_17
timestamp 1764626446
transform -1 0 668 0 1 20108
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_18
timestamp 1764626446
transform -1 0 668 0 1 22532
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_19
timestamp 1764626446
transform -1 0 668 0 1 23744
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_20
timestamp 1764626446
transform -1 0 668 0 1 24956
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_21
timestamp 1764626446
transform -1 0 668 0 1 26168
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_22
timestamp 1764626446
transform -1 0 668 0 1 27380
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_23
timestamp 1764626446
transform -1 0 668 0 1 28592
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_24
timestamp 1764626446
transform -1 0 668 0 1 29804
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_25
timestamp 1764626446
transform -1 0 668 0 1 31016
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_26
timestamp 1764626446
transform -1 0 668 0 1 32228
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_27
timestamp 1764626446
transform -1 0 668 0 1 33440
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_28
timestamp 1764626446
transform -1 0 668 0 1 34652
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_29
timestamp 1764626446
transform -1 0 668 0 1 35864
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_30
timestamp 1764626446
transform -1 0 668 0 1 37076
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_31
timestamp 1764626446
transform -1 0 668 0 1 1928
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_32
timestamp 1764626446
transform -1 0 668 0 -1 38540
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_33
timestamp 1764626446
transform -1 0 668 0 -1 37328
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_34
timestamp 1764626446
transform -1 0 668 0 -1 36116
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_35
timestamp 1764626446
transform -1 0 668 0 -1 34904
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_36
timestamp 1764626446
transform -1 0 668 0 -1 33692
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_37
timestamp 1764626446
transform -1 0 668 0 -1 32480
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_38
timestamp 1764626446
transform -1 0 668 0 -1 31268
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_39
timestamp 1764626446
transform -1 0 668 0 -1 30056
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_40
timestamp 1764626446
transform -1 0 668 0 -1 28844
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_41
timestamp 1764626446
transform -1 0 668 0 -1 27632
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_42
timestamp 1764626446
transform -1 0 668 0 -1 26420
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_43
timestamp 1764626446
transform -1 0 668 0 -1 25208
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_44
timestamp 1764626446
transform -1 0 668 0 -1 23996
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_45
timestamp 1764626446
transform -1 0 668 0 -1 22784
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_46
timestamp 1764626446
transform -1 0 668 0 -1 20360
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_47
timestamp 1764626446
transform -1 0 668 0 -1 21572
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_48
timestamp 1764626446
transform -1 0 668 0 -1 19148
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_49
timestamp 1764626446
transform -1 0 668 0 -1 17936
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_50
timestamp 1764626446
transform -1 0 668 0 -1 16724
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_51
timestamp 1764626446
transform -1 0 668 0 -1 15512
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_52
timestamp 1764626446
transform -1 0 668 0 -1 14300
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_53
timestamp 1764626446
transform -1 0 668 0 -1 13088
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_54
timestamp 1764626446
transform -1 0 668 0 -1 11876
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_55
timestamp 1764626446
transform -1 0 668 0 -1 10664
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_56
timestamp 1764626446
transform -1 0 668 0 -1 9452
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_57
timestamp 1764626446
transform -1 0 668 0 -1 8240
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_58
timestamp 1764626446
transform -1 0 668 0 -1 7028
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_59
timestamp 1764626446
transform -1 0 668 0 -1 5816
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_60
timestamp 1764626446
transform -1 0 668 0 -1 4604
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_61
timestamp 1764626446
transform -1 0 668 0 -1 3392
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_62
timestamp 1764626446
transform -1 0 668 0 -1 968
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_63
timestamp 1764626446
transform -1 0 668 0 -1 2180
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_64
timestamp 1764626446
transform -1 0 668 0 1 39500
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_65
timestamp 1764626446
transform -1 0 668 0 -1 39752
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_66
timestamp 1764626446
transform -1 0 668 0 1 40712
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_67
timestamp 1764626446
transform -1 0 668 0 -1 40964
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_68
timestamp 1764626446
transform -1 0 668 0 1 41924
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_69
timestamp 1764626446
transform -1 0 668 0 -1 42176
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_70
timestamp 1764626446
transform -1 0 668 0 1 43136
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_71
timestamp 1764626446
transform -1 0 668 0 -1 43388
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_72
timestamp 1764626446
transform -1 0 668 0 1 44348
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_73
timestamp 1764626446
transform -1 0 668 0 -1 44600
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_74
timestamp 1764626446
transform -1 0 668 0 1 45560
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_75
timestamp 1764626446
transform -1 0 668 0 -1 45812
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_76
timestamp 1764626446
transform -1 0 668 0 1 46772
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_77
timestamp 1764626446
transform -1 0 668 0 -1 47024
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_78
timestamp 1764626446
transform -1 0 668 0 1 47984
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_79
timestamp 1764626446
transform -1 0 668 0 -1 48236
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_80
timestamp 1764626446
transform -1 0 668 0 1 49196
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_81
timestamp 1764626446
transform -1 0 668 0 -1 49448
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_82
timestamp 1764626446
transform -1 0 668 0 1 50408
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_83
timestamp 1764626446
transform -1 0 668 0 -1 50660
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_84
timestamp 1764626446
transform -1 0 668 0 1 51620
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_85
timestamp 1764626446
transform -1 0 668 0 -1 51872
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_86
timestamp 1764626446
transform -1 0 668 0 1 52832
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_87
timestamp 1764626446
transform -1 0 668 0 -1 53084
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_88
timestamp 1764626446
transform -1 0 668 0 1 54044
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_89
timestamp 1764626446
transform -1 0 668 0 -1 54296
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_90
timestamp 1764626446
transform -1 0 668 0 1 55256
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_91
timestamp 1764626446
transform -1 0 668 0 -1 55508
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_92
timestamp 1764626446
transform -1 0 668 0 1 56468
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_93
timestamp 1764626446
transform -1 0 668 0 -1 56720
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_94
timestamp 1764626446
transform -1 0 668 0 1 57680
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_95
timestamp 1764626446
transform -1 0 668 0 -1 57932
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_96
timestamp 1764626446
transform -1 0 668 0 1 58892
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_97
timestamp 1764626446
transform -1 0 668 0 -1 59144
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_98
timestamp 1764626446
transform -1 0 668 0 1 60104
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_99
timestamp 1764626446
transform -1 0 668 0 -1 60356
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_100
timestamp 1764626446
transform -1 0 668 0 1 61316
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_101
timestamp 1764626446
transform -1 0 668 0 -1 61568
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_102
timestamp 1764626446
transform -1 0 668 0 1 62528
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_103
timestamp 1764626446
transform -1 0 668 0 -1 62780
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_104
timestamp 1764626446
transform -1 0 668 0 1 63740
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_105
timestamp 1764626446
transform -1 0 668 0 -1 63992
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_106
timestamp 1764626446
transform -1 0 668 0 1 64952
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_107
timestamp 1764626446
transform -1 0 668 0 -1 65204
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_108
timestamp 1764626446
transform -1 0 668 0 1 66164
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_109
timestamp 1764626446
transform -1 0 668 0 -1 66416
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_110
timestamp 1764626446
transform -1 0 668 0 1 67376
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_111
timestamp 1764626446
transform -1 0 668 0 -1 67628
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_112
timestamp 1764626446
transform -1 0 668 0 1 68588
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_113
timestamp 1764626446
transform -1 0 668 0 -1 68840
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_114
timestamp 1764626446
transform -1 0 668 0 1 69800
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_115
timestamp 1764626446
transform -1 0 668 0 -1 70052
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_116
timestamp 1764626446
transform -1 0 668 0 1 71012
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_117
timestamp 1764626446
transform -1 0 668 0 -1 71264
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_118
timestamp 1764626446
transform -1 0 668 0 1 72224
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_119
timestamp 1764626446
transform -1 0 668 0 -1 72476
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_120
timestamp 1764626446
transform -1 0 668 0 1 73436
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_121
timestamp 1764626446
transform -1 0 668 0 -1 73688
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_122
timestamp 1764626446
transform -1 0 668 0 1 74648
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_123
timestamp 1764626446
transform -1 0 668 0 -1 74900
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_124
timestamp 1764626446
transform -1 0 668 0 1 75860
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_125
timestamp 1764626446
transform -1 0 668 0 -1 76112
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_126
timestamp 1764626446
transform -1 0 668 0 1 77072
box 30 89 570 797
use 018SRAM_cell1_cutPC_3v1024x8m81  018SRAM_cell1_cutPC_3v1024x8m81_127
timestamp 1764626446
transform -1 0 668 0 -1 77324
box 30 89 570 797
<< labels >>
rlabel metal1 s 572 19623 572 19623 4 VDD
rlabel metal1 s 570 20097 570 20097 4 VSS
rlabel metal1 s 570 983 570 983 4 VSS
rlabel metal1 s 567 232 567 232 4 VDD
<< end >>
