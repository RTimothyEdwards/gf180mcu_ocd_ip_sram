magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< psubdiff >>
rect -571 23 571 55
rect -571 -23 -537 23
rect 537 -23 571 23
rect -571 -56 571 -23
<< psubdiffcont >>
rect -537 -23 537 23
<< metal1 >>
rect -565 23 565 49
rect -565 -23 -537 23
rect 537 -23 565 23
rect -565 -49 565 -23
<< end >>
