magic
tech gf180mcuD
magscale 1 10
timestamp 1764700137
<< metal2 >>
rect -561 28 562 46
rect -561 -28 -545 28
rect 545 -28 562 28
rect -561 -46 562 -28
<< via2 >>
rect -545 -28 545 28
<< metal3 >>
rect -562 28 562 46
rect -562 -28 -545 28
rect 545 -28 562 28
rect -562 -46 562 -28
<< end >>
