magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< polysilicon >>
rect -14 211 41 245
rect -14 -34 41 0
use nmos_5p04310591302010_256x8m81  nmos_5p04310591302010_256x8m81_0
timestamp 1763766357
transform 1 0 -14 0 1 0
box -88 -44 144 255
<< end >>
