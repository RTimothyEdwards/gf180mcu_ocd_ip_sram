VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_ocd_ip_sram__sram256x8m8wm1
  CLASS BLOCK ;
  FOREIGN gf180mcu_ocd_ip_sram__sram256x8m8wm1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 301.300 BY 224.930 ;
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 103.965 0.700 104.750 6.000 ;
        RECT 103.960 0.000 104.750 0.700 ;
    END
  END A[7]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 188.200 0.000 188.985 6.000 ;
    END
  END A[6]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 190.455 0.000 191.240 6.000 ;
    END
  END A[5]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 193.070 0.000 193.855 6.000 ;
    END
  END A[4]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 196.925 0.000 197.710 6.000 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 108.005 0.000 108.790 6.000 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 113.930 0.000 114.715 6.000 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 119.850 0.000 120.630 6.000 ;
    END
  END A[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 176.195 0.000 176.980 6.000 ;
    END
  END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.738400 ;
    PORT
      LAYER Metal2 ;
        RECT 97.775 0.000 98.560 6.000 ;
    END
  END CLK
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 291.200 5.030 291.985 6.000 ;
        RECT 290.800 4.305 291.985 5.030 ;
        RECT 290.800 0.000 291.585 4.305 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 254.645 4.245 254.930 6.000 ;
        RECT 254.605 0.000 255.385 4.245 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 249.530 4.245 249.810 6.000 ;
        RECT 249.235 0.000 250.020 4.245 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 212.255 4.355 212.625 6.000 ;
        RECT 212.255 4.350 213.940 4.355 ;
        RECT 212.255 3.985 214.845 4.350 ;
        RECT 214.060 0.000 214.845 3.985 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 85.695 4.850 86.000 6.000 ;
        RECT 83.280 4.545 86.000 4.850 ;
        RECT 83.280 0.000 84.065 4.545 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 48.730 5.425 49.015 6.000 ;
        RECT 47.595 5.140 49.015 5.425 ;
        RECT 47.595 4.160 47.880 5.140 ;
        RECT 47.085 3.720 47.880 4.160 ;
        RECT 47.085 0.000 47.870 3.720 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 43.215 5.290 43.540 6.000 ;
        RECT 43.180 4.170 43.540 5.290 ;
        RECT 42.720 0.000 43.505 4.170 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 6.520 0.000 7.305 6.000 ;
    END
  END D[0]
  PIN GWEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.141600 ;
    PORT
      LAYER Metal2 ;
        RECT 142.055 0.000 142.840 6.000 ;
    END
  END GWEN
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 285.870 4.245 286.200 6.000 ;
        RECT 285.490 0.000 286.275 4.245 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 257.025 4.245 257.345 6.000 ;
        RECT 256.960 0.000 257.740 4.245 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 247.175 4.245 247.460 6.000 ;
        RECT 246.880 0.000 247.665 4.245 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 217.860 4.705 218.190 6.000 ;
        RECT 217.860 4.695 220.060 4.705 ;
        RECT 217.860 4.375 220.135 4.695 ;
        RECT 219.350 0.000 220.135 4.375 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 77.980 4.130 78.315 6.000 ;
        RECT 77.975 0.000 78.760 4.130 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 51.250 5.450 51.580 6.000 ;
        RECT 49.960 5.120 51.580 5.450 ;
        RECT 49.960 4.160 50.290 5.120 ;
        RECT 49.440 3.710 50.290 4.160 ;
        RECT 49.440 0.000 50.225 3.710 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 41.545 4.725 41.875 6.000 ;
        RECT 40.840 4.395 41.875 4.725 ;
        RECT 40.840 4.200 41.170 4.395 ;
        RECT 40.365 3.555 41.170 4.200 ;
        RECT 40.365 0.000 41.145 3.555 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 12.255 5.780 12.585 6.000 ;
        RECT 12.255 5.450 14.415 5.780 ;
        RECT 14.085 4.245 14.415 5.450 ;
        RECT 13.830 0.000 14.610 4.245 ;
    END
  END Q[0]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT 103.900 218.930 194.020 219.810 ;
        RECT 7.680 5.780 25.360 6.000 ;
        RECT 29.080 5.780 64.190 6.000 ;
        RECT 29.080 5.770 46.760 5.780 ;
        RECT 67.910 5.770 85.590 6.000 ;
        RECT 212.985 5.780 230.665 6.000 ;
        RECT 234.385 5.785 269.745 6.000 ;
        RECT 234.385 5.770 252.065 5.785 ;
        RECT 273.465 5.775 291.145 6.000 ;
      LAYER Metal1 ;
        RECT 4.845 214.375 5.975 215.090 ;
        RECT 4.845 213.675 6.000 214.375 ;
        RECT 295.440 214.170 296.570 215.175 ;
        RECT 295.300 213.790 296.570 214.170 ;
        RECT 4.845 212.660 5.975 213.675 ;
        RECT 295.440 212.745 296.570 213.790 ;
        RECT 4.845 208.315 5.975 209.030 ;
        RECT 4.845 207.615 6.000 208.315 ;
        RECT 295.440 208.110 296.570 209.115 ;
        RECT 295.300 207.730 296.570 208.110 ;
        RECT 4.845 206.600 5.975 207.615 ;
        RECT 295.440 206.685 296.570 207.730 ;
        RECT 4.845 202.255 5.975 202.970 ;
        RECT 4.845 201.555 6.000 202.255 ;
        RECT 295.440 202.050 296.570 203.055 ;
        RECT 295.300 201.670 296.570 202.050 ;
        RECT 4.845 200.540 5.975 201.555 ;
        RECT 295.440 200.625 296.570 201.670 ;
        RECT 4.845 196.195 5.975 196.910 ;
        RECT 4.845 195.495 6.000 196.195 ;
        RECT 295.440 195.990 296.570 196.995 ;
        RECT 295.300 195.610 296.570 195.990 ;
        RECT 4.845 194.480 5.975 195.495 ;
        RECT 295.440 194.565 296.570 195.610 ;
        RECT 4.845 190.135 5.975 190.850 ;
        RECT 4.845 189.435 6.000 190.135 ;
        RECT 295.440 189.930 296.570 190.935 ;
        RECT 295.300 189.550 296.570 189.930 ;
        RECT 4.845 188.420 5.975 189.435 ;
        RECT 295.440 188.505 296.570 189.550 ;
        RECT 4.845 184.075 5.975 184.790 ;
        RECT 4.845 183.375 6.000 184.075 ;
        RECT 295.440 183.870 296.570 184.875 ;
        RECT 295.300 183.490 296.570 183.870 ;
        RECT 4.845 182.360 5.975 183.375 ;
        RECT 295.440 182.445 296.570 183.490 ;
        RECT 4.845 178.015 5.975 178.730 ;
        RECT 4.845 177.315 6.000 178.015 ;
        RECT 295.440 177.810 296.570 178.815 ;
        RECT 295.300 177.430 296.570 177.810 ;
        RECT 4.845 176.300 5.975 177.315 ;
        RECT 295.440 176.385 296.570 177.430 ;
        RECT 4.845 171.955 5.975 172.670 ;
        RECT 4.845 171.255 6.000 171.955 ;
        RECT 295.440 171.750 296.570 172.755 ;
        RECT 295.300 171.370 296.570 171.750 ;
        RECT 4.845 170.240 5.975 171.255 ;
        RECT 295.440 170.325 296.570 171.370 ;
        RECT 4.845 165.895 5.975 166.610 ;
        RECT 4.845 165.195 6.000 165.895 ;
        RECT 295.440 165.690 296.570 166.695 ;
        RECT 295.300 165.310 296.570 165.690 ;
        RECT 4.845 164.180 5.975 165.195 ;
        RECT 295.440 164.265 296.570 165.310 ;
        RECT 4.845 159.835 5.975 160.550 ;
        RECT 4.845 159.135 6.000 159.835 ;
        RECT 295.440 159.630 296.570 160.635 ;
        RECT 295.300 159.250 296.570 159.630 ;
        RECT 4.845 158.120 5.975 159.135 ;
        RECT 295.440 158.205 296.570 159.250 ;
        RECT 4.845 153.775 5.975 154.490 ;
        RECT 4.845 153.075 6.000 153.775 ;
        RECT 295.440 153.570 296.570 154.575 ;
        RECT 295.300 153.190 296.570 153.570 ;
        RECT 4.845 152.060 5.975 153.075 ;
        RECT 295.440 152.145 296.570 153.190 ;
        RECT 4.845 147.715 5.975 148.430 ;
        RECT 4.845 147.015 6.000 147.715 ;
        RECT 295.440 147.510 296.570 148.515 ;
        RECT 295.300 147.130 296.570 147.510 ;
        RECT 4.845 146.000 5.975 147.015 ;
        RECT 295.440 146.085 296.570 147.130 ;
        RECT 4.845 141.655 5.975 142.370 ;
        RECT 4.845 140.955 6.000 141.655 ;
        RECT 295.440 141.450 296.570 142.455 ;
        RECT 295.300 141.070 296.570 141.450 ;
        RECT 4.845 139.940 5.975 140.955 ;
        RECT 295.440 140.025 296.570 141.070 ;
        RECT 4.845 135.595 5.975 136.310 ;
        RECT 4.845 134.895 6.000 135.595 ;
        RECT 295.440 135.390 296.570 136.395 ;
        RECT 295.300 135.010 296.570 135.390 ;
        RECT 4.845 133.880 5.975 134.895 ;
        RECT 295.440 133.965 296.570 135.010 ;
        RECT 4.845 129.535 5.975 130.250 ;
        RECT 4.845 128.835 6.000 129.535 ;
        RECT 295.440 129.330 296.570 130.335 ;
        RECT 295.300 128.950 296.570 129.330 ;
        RECT 4.845 127.820 5.975 128.835 ;
        RECT 295.440 127.905 296.570 128.950 ;
        RECT 4.845 123.475 5.975 124.190 ;
        RECT 4.845 122.775 6.000 123.475 ;
        RECT 295.440 123.270 296.570 124.275 ;
        RECT 295.300 122.890 296.570 123.270 ;
        RECT 4.845 121.760 5.975 122.775 ;
        RECT 295.440 121.845 296.570 122.890 ;
        RECT 4.845 117.415 5.975 118.130 ;
        RECT 4.845 116.715 6.000 117.415 ;
        RECT 295.440 117.210 296.570 118.215 ;
        RECT 295.300 116.830 296.570 117.210 ;
        RECT 4.845 115.700 5.975 116.715 ;
        RECT 295.440 115.785 296.570 116.830 ;
        RECT 93.700 5.990 95.245 6.000 ;
      LAYER Metal2 ;
        RECT 2.470 221.980 298.830 222.130 ;
        RECT 2.465 218.930 298.830 221.980 ;
        RECT 2.465 218.630 6.000 218.930 ;
        RECT 295.300 218.630 298.830 218.930 ;
        RECT 2.465 215.090 5.970 218.630 ;
        RECT 295.445 215.310 298.830 218.630 ;
        RECT 2.465 212.660 5.975 215.090 ;
        RECT 2.465 209.030 5.970 212.660 ;
        RECT 2.465 206.600 5.975 209.030 ;
        RECT 2.465 202.970 5.970 206.600 ;
        RECT 2.465 200.540 5.975 202.970 ;
        RECT 2.465 196.910 5.970 200.540 ;
        RECT 2.465 194.480 5.975 196.910 ;
        RECT 2.465 190.850 5.970 194.480 ;
        RECT 2.465 188.420 5.975 190.850 ;
        RECT 2.465 184.790 5.970 188.420 ;
        RECT 2.465 182.360 5.975 184.790 ;
        RECT 2.465 178.730 5.970 182.360 ;
        RECT 2.465 176.300 5.975 178.730 ;
        RECT 2.465 172.670 5.970 176.300 ;
        RECT 2.465 170.240 5.975 172.670 ;
        RECT 2.465 166.610 5.970 170.240 ;
        RECT 295.440 168.360 298.830 215.310 ;
        RECT 2.465 164.180 5.975 166.610 ;
        RECT 2.465 160.550 5.970 164.180 ;
        RECT 2.465 158.120 5.975 160.550 ;
        RECT 2.465 154.490 5.970 158.120 ;
        RECT 2.465 152.060 5.975 154.490 ;
        RECT 2.465 148.430 5.970 152.060 ;
        RECT 2.465 146.000 5.975 148.430 ;
        RECT 2.465 142.370 5.970 146.000 ;
        RECT 2.465 139.940 5.975 142.370 ;
        RECT 2.465 136.310 5.970 139.940 ;
        RECT 2.465 133.880 5.975 136.310 ;
        RECT 2.465 130.250 5.970 133.880 ;
        RECT 2.465 127.820 5.975 130.250 ;
        RECT 2.465 124.190 5.970 127.820 ;
        RECT 2.465 121.760 5.975 124.190 ;
        RECT 2.465 118.130 5.970 121.760 ;
        RECT 2.465 115.700 5.975 118.130 ;
        RECT 2.465 110.435 5.970 115.700 ;
        RECT 295.440 110.435 298.835 168.360 ;
        RECT 2.465 4.330 5.975 110.435 ;
        RECT 26.795 4.830 27.580 6.000 ;
        RECT 65.605 4.830 66.390 6.000 ;
        RECT 2.465 1.410 5.970 4.330 ;
        RECT 88.750 4.285 89.535 6.000 ;
        RECT 93.695 5.965 95.245 6.000 ;
        RECT 131.250 5.180 132.035 6.000 ;
        RECT 137.620 5.180 138.405 6.000 ;
        RECT 207.850 4.315 208.635 6.000 ;
        RECT 232.070 4.830 232.855 6.000 ;
        RECT 271.220 4.810 272.005 6.000 ;
        RECT 295.330 4.330 298.835 110.435 ;
        RECT 2.470 0.985 5.970 1.410 ;
        RECT 295.330 0.985 298.830 4.330 ;
      LAYER Metal3 ;
        RECT 5.090 222.130 8.585 224.930 ;
        RECT 14.480 222.130 17.975 224.930 ;
        RECT 24.630 222.130 28.125 224.930 ;
        RECT 33.380 222.130 36.875 224.930 ;
        RECT 44.170 222.130 47.665 224.930 ;
        RECT 52.280 222.130 55.775 224.930 ;
        RECT 63.710 222.130 67.205 224.930 ;
        RECT 72.285 222.130 75.780 224.930 ;
        RECT 84.685 222.130 88.180 224.930 ;
        RECT 93.000 222.130 96.495 224.930 ;
        RECT 107.485 222.130 110.980 224.930 ;
        RECT 123.950 222.130 127.445 224.930 ;
        RECT 135.045 222.130 138.540 224.930 ;
        RECT 144.305 222.130 147.800 224.930 ;
        RECT 157.740 222.130 161.235 224.930 ;
        RECT 162.095 222.130 165.590 224.930 ;
        RECT 171.155 222.130 174.650 224.930 ;
        RECT 183.990 222.130 187.485 224.930 ;
        RECT 189.915 222.130 193.410 224.930 ;
        RECT 201.415 222.130 204.910 224.930 ;
        RECT 210.520 222.130 214.015 224.930 ;
        RECT 221.995 222.130 225.490 224.930 ;
        RECT 230.060 222.130 233.555 224.930 ;
        RECT 240.895 222.130 244.390 224.930 ;
        RECT 249.600 222.130 253.095 224.930 ;
        RECT 259.795 222.130 263.290 224.930 ;
        RECT 269.140 222.130 272.635 224.930 ;
        RECT 279.300 222.130 282.795 224.930 ;
        RECT 290.115 222.130 293.610 224.930 ;
        RECT 295.330 222.130 298.825 224.930 ;
        RECT 0.000 218.930 301.300 222.130 ;
        RECT 0.000 218.630 6.000 218.930 ;
        RECT 295.300 218.630 301.300 218.930 ;
        RECT 5.090 218.625 6.000 218.630 ;
        RECT 296.440 215.175 301.300 215.185 ;
        RECT 0.000 212.650 5.975 215.100 ;
        RECT 295.440 212.745 301.300 215.175 ;
        RECT 296.440 212.735 301.300 212.745 ;
        RECT 296.440 209.115 301.300 209.125 ;
        RECT 0.000 206.590 5.975 209.040 ;
        RECT 295.440 206.685 301.300 209.115 ;
        RECT 296.440 206.675 301.300 206.685 ;
        RECT 296.440 203.055 301.300 203.065 ;
        RECT 0.000 200.530 5.975 202.980 ;
        RECT 295.440 200.625 301.300 203.055 ;
        RECT 296.440 200.615 301.300 200.625 ;
        RECT 296.440 196.995 301.300 197.005 ;
        RECT 0.000 194.470 5.975 196.920 ;
        RECT 295.440 194.565 301.300 196.995 ;
        RECT 296.440 194.555 301.300 194.565 ;
        RECT 296.440 190.935 301.300 190.945 ;
        RECT 0.000 188.410 5.975 190.860 ;
        RECT 295.440 188.505 301.300 190.935 ;
        RECT 296.440 188.495 301.300 188.505 ;
        RECT 296.440 184.875 301.300 184.885 ;
        RECT 0.000 182.350 5.975 184.800 ;
        RECT 295.440 182.445 301.300 184.875 ;
        RECT 296.440 182.435 301.300 182.445 ;
        RECT 296.440 178.815 301.300 178.825 ;
        RECT 0.000 176.290 5.975 178.740 ;
        RECT 295.440 176.385 301.300 178.815 ;
        RECT 296.440 176.375 301.300 176.385 ;
        RECT 296.440 172.755 301.300 172.765 ;
        RECT 0.000 170.230 5.975 172.680 ;
        RECT 295.440 170.325 301.300 172.755 ;
        RECT 296.440 170.315 301.300 170.325 ;
        RECT 296.440 166.695 301.300 166.705 ;
        RECT 0.000 164.170 5.975 166.620 ;
        RECT 295.440 164.265 301.300 166.695 ;
        RECT 296.440 164.255 301.300 164.265 ;
        RECT 296.440 160.635 301.300 160.645 ;
        RECT 0.000 158.110 5.975 160.560 ;
        RECT 295.440 158.205 301.300 160.635 ;
        RECT 296.440 158.195 301.300 158.205 ;
        RECT 296.440 154.575 301.300 154.585 ;
        RECT 0.000 152.050 5.975 154.500 ;
        RECT 295.440 152.145 301.300 154.575 ;
        RECT 296.440 152.135 301.300 152.145 ;
        RECT 296.440 148.515 301.300 148.525 ;
        RECT 0.000 145.990 5.975 148.440 ;
        RECT 295.440 146.085 301.300 148.515 ;
        RECT 296.440 146.075 301.300 146.085 ;
        RECT 296.440 142.455 301.300 142.465 ;
        RECT 0.000 139.930 5.975 142.380 ;
        RECT 295.440 140.025 301.300 142.455 ;
        RECT 296.440 140.015 301.300 140.025 ;
        RECT 296.440 136.395 301.300 136.405 ;
        RECT 0.000 133.870 5.975 136.320 ;
        RECT 295.440 133.965 301.300 136.395 ;
        RECT 296.440 133.955 301.300 133.965 ;
        RECT 296.440 130.335 301.300 130.345 ;
        RECT 0.000 127.810 5.975 130.260 ;
        RECT 295.440 127.905 301.300 130.335 ;
        RECT 296.440 127.895 301.300 127.905 ;
        RECT 296.440 124.275 301.300 124.285 ;
        RECT 0.000 121.750 5.975 124.200 ;
        RECT 295.440 121.845 301.300 124.275 ;
        RECT 296.440 121.835 301.300 121.845 ;
        RECT 296.440 118.215 301.300 118.225 ;
        RECT 0.000 115.690 5.975 118.140 ;
        RECT 295.440 115.785 301.300 118.215 ;
        RECT 296.440 115.775 301.300 115.785 ;
        RECT 0.000 109.905 3.545 109.910 ;
        RECT 297.750 109.905 301.300 109.910 ;
        RECT 0.000 102.880 6.000 109.905 ;
        RECT 295.300 102.880 301.300 109.905 ;
        RECT 0.000 96.170 5.975 102.880 ;
        RECT 295.335 96.170 301.300 102.880 ;
        RECT 0.000 95.175 6.000 96.170 ;
        RECT 295.300 95.175 301.300 96.170 ;
        RECT 300.600 95.170 301.300 95.175 ;
        RECT 0.000 78.350 3.545 78.355 ;
        RECT 297.750 78.350 301.300 78.355 ;
        RECT 0.000 76.400 5.975 78.350 ;
        RECT 295.335 76.400 301.300 78.350 ;
        RECT 0.000 74.855 6.000 76.400 ;
        RECT 0.010 74.850 6.000 74.855 ;
        RECT 295.300 74.850 301.300 76.400 ;
        RECT 297.750 67.740 301.300 67.750 ;
        RECT 0.010 67.735 6.000 67.740 ;
        RECT 0.000 58.210 6.000 67.735 ;
        RECT 295.300 58.210 301.300 67.740 ;
        RECT 0.000 58.205 0.700 58.210 ;
        RECT 300.600 58.205 301.300 58.210 ;
        RECT 0.000 47.315 3.545 47.325 ;
        RECT 300.600 47.315 301.300 47.320 ;
        RECT 0.000 44.810 6.000 47.315 ;
        RECT 295.300 44.810 301.300 47.315 ;
        RECT 0.000 42.955 5.975 44.810 ;
        RECT 295.335 42.970 301.300 44.810 ;
        RECT 0.000 40.125 6.000 42.955 ;
        RECT 0.010 40.120 6.000 40.125 ;
        RECT 295.300 40.120 301.300 42.970 ;
        RECT 0.010 40.020 5.975 40.120 ;
        RECT 295.335 40.020 301.300 40.120 ;
        RECT 297.750 40.010 301.300 40.020 ;
        RECT 0.000 31.295 3.545 31.300 ;
        RECT 295.300 31.295 295.365 31.325 ;
        RECT 300.600 31.295 301.300 31.300 ;
        RECT 0.000 26.530 6.000 31.295 ;
        RECT 0.010 26.525 6.000 26.530 ;
        RECT 295.300 26.525 301.300 31.295 ;
        RECT 0.000 19.345 3.545 19.350 ;
        RECT 297.750 19.345 301.300 19.350 ;
        RECT 0.000 17.750 6.000 19.345 ;
        RECT 0.000 15.795 5.995 17.750 ;
        RECT 295.300 17.745 301.300 19.345 ;
        RECT 295.315 15.805 301.300 17.745 ;
        RECT 0.000 14.210 6.000 15.795 ;
        RECT 0.010 14.205 6.000 14.210 ;
        RECT 295.300 14.205 301.300 15.805 ;
        RECT 0.000 6.000 6.000 7.810 ;
        RECT 295.300 6.000 301.300 7.810 ;
        RECT 0.000 4.310 301.300 6.000 ;
        RECT 0.000 4.290 0.700 4.310 ;
        RECT 2.465 0.000 5.970 4.310 ;
        RECT 7.135 0.000 10.635 4.310 ;
        RECT 12.045 0.000 15.545 4.310 ;
        RECT 20.445 0.000 23.945 4.310 ;
        RECT 24.645 0.000 28.145 4.310 ;
        RECT 28.845 0.000 32.345 4.310 ;
        RECT 37.245 0.000 40.745 4.310 ;
        RECT 43.550 0.000 47.050 4.310 ;
        RECT 49.845 0.000 53.345 4.310 ;
        RECT 58.245 0.000 61.745 4.310 ;
        RECT 62.445 0.000 65.945 4.310 ;
        RECT 66.645 0.000 70.145 4.310 ;
        RECT 76.685 0.000 80.185 4.310 ;
        RECT 80.885 0.000 84.385 4.310 ;
        RECT 85.435 0.000 88.935 4.310 ;
        RECT 89.985 0.000 93.485 4.310 ;
        RECT 94.535 0.000 98.035 4.310 ;
        RECT 99.085 0.000 102.585 4.310 ;
        RECT 103.635 0.000 107.135 4.310 ;
        RECT 126.105 0.000 129.605 4.310 ;
        RECT 137.295 0.000 140.795 4.310 ;
        RECT 148.515 0.000 152.015 4.310 ;
        RECT 156.915 0.000 160.415 4.310 ;
        RECT 165.315 0.000 168.815 4.310 ;
        RECT 169.980 0.000 173.480 4.310 ;
        RECT 174.565 0.000 178.065 4.310 ;
        RECT 190.600 0.000 194.100 4.310 ;
        RECT 195.150 0.000 198.650 4.310 ;
        RECT 199.700 4.205 221.530 4.310 ;
        RECT 199.700 0.000 203.200 4.205 ;
        RECT 204.250 0.000 207.750 4.205 ;
        RECT 208.800 0.000 212.300 4.205 ;
        RECT 213.350 0.000 216.850 4.205 ;
        RECT 218.030 0.000 221.530 4.205 ;
        RECT 227.960 0.000 231.460 4.310 ;
        RECT 232.160 0.000 235.660 4.310 ;
        RECT 236.360 0.000 239.860 4.310 ;
        RECT 244.760 0.000 248.260 4.310 ;
        RECT 251.055 0.000 254.555 4.310 ;
        RECT 257.360 0.000 260.860 4.310 ;
        RECT 265.760 0.000 269.260 4.310 ;
        RECT 269.960 0.000 273.460 4.310 ;
        RECT 274.160 0.000 277.660 4.310 ;
        RECT 283.560 0.000 287.060 4.310 ;
        RECT 288.465 0.000 291.965 4.310 ;
        RECT 295.330 0.000 298.830 4.310 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.985 220.405 300.315 223.940 ;
        RECT 0.985 218.075 4.485 220.405 ;
        RECT 7.150 218.930 7.970 220.405 ;
        RECT 26.690 218.930 27.510 220.405 ;
        RECT 46.230 218.930 47.050 220.405 ;
        RECT 65.770 218.930 66.590 220.405 ;
        RECT 85.300 218.930 86.120 220.405 ;
        RECT 90.140 218.930 92.685 220.405 ;
        RECT 96.620 220.070 102.185 220.405 ;
        RECT 95.855 218.930 102.185 220.070 ;
        RECT 119.790 218.930 122.545 220.405 ;
        RECT 140.215 218.930 142.065 220.405 ;
        RECT 153.080 218.930 155.970 220.405 ;
        RECT 175.340 218.930 178.195 220.405 ;
        RECT 194.845 218.930 202.075 220.405 ;
        RECT 204.765 218.930 207.310 220.405 ;
        RECT 212.580 218.930 213.400 220.405 ;
        RECT 232.120 218.930 232.940 220.405 ;
        RECT 251.660 218.930 252.480 220.405 ;
        RECT 271.200 218.930 272.020 220.405 ;
        RECT 290.730 218.930 291.550 220.405 ;
        RECT 0.985 217.925 4.490 218.075 ;
        RECT 0.985 216.120 6.000 217.925 ;
        RECT 0.985 212.825 4.490 216.120 ;
        RECT 0.985 212.015 4.485 212.825 ;
        RECT 0.985 211.865 4.490 212.015 ;
        RECT 0.985 210.060 6.000 211.865 ;
        RECT 0.985 206.765 4.490 210.060 ;
        RECT 0.985 205.955 4.485 206.765 ;
        RECT 0.985 205.805 4.490 205.955 ;
        RECT 0.985 204.000 6.000 205.805 ;
        RECT 0.985 200.705 4.490 204.000 ;
        RECT 0.985 199.895 4.485 200.705 ;
        RECT 0.985 199.745 4.490 199.895 ;
        RECT 0.985 197.940 6.000 199.745 ;
        RECT 0.985 194.645 4.490 197.940 ;
        RECT 0.985 193.835 4.485 194.645 ;
        RECT 0.985 193.685 4.490 193.835 ;
        RECT 0.985 191.880 6.000 193.685 ;
        RECT 0.985 188.585 4.490 191.880 ;
        RECT 0.985 187.775 4.485 188.585 ;
        RECT 0.985 187.625 4.490 187.775 ;
        RECT 0.985 185.820 6.000 187.625 ;
        RECT 0.985 182.525 4.490 185.820 ;
        RECT 0.985 181.715 4.485 182.525 ;
        RECT 0.985 181.565 4.490 181.715 ;
        RECT 0.985 179.760 6.000 181.565 ;
        RECT 0.985 176.465 4.490 179.760 ;
        RECT 0.985 175.655 4.485 176.465 ;
        RECT 0.985 175.505 4.490 175.655 ;
        RECT 0.985 173.700 6.000 175.505 ;
        RECT 0.985 170.405 4.490 173.700 ;
        RECT 0.985 169.595 4.485 170.405 ;
        RECT 0.985 169.445 4.490 169.595 ;
        RECT 0.985 167.640 6.000 169.445 ;
        RECT 0.985 164.345 4.490 167.640 ;
        RECT 0.985 163.535 4.485 164.345 ;
        RECT 0.985 163.385 4.490 163.535 ;
        RECT 0.985 161.580 6.000 163.385 ;
        RECT 0.985 158.285 4.490 161.580 ;
        RECT 0.985 157.475 4.485 158.285 ;
        RECT 0.985 157.325 4.490 157.475 ;
        RECT 0.985 155.520 6.000 157.325 ;
        RECT 0.985 152.225 4.490 155.520 ;
        RECT 0.985 151.415 4.485 152.225 ;
        RECT 0.985 151.265 4.490 151.415 ;
        RECT 0.985 149.460 6.000 151.265 ;
        RECT 0.985 146.165 4.490 149.460 ;
        RECT 0.985 145.355 4.485 146.165 ;
        RECT 0.985 145.205 4.490 145.355 ;
        RECT 0.985 143.400 6.000 145.205 ;
        RECT 0.985 140.105 4.490 143.400 ;
        RECT 0.985 139.295 4.485 140.105 ;
        RECT 0.985 139.145 4.490 139.295 ;
        RECT 0.985 137.340 6.000 139.145 ;
        RECT 0.985 134.045 4.490 137.340 ;
        RECT 0.985 133.235 4.485 134.045 ;
        RECT 0.985 133.085 4.490 133.235 ;
        RECT 0.985 131.280 6.000 133.085 ;
        RECT 0.985 127.985 4.490 131.280 ;
        RECT 0.985 127.175 4.485 127.985 ;
        RECT 0.985 127.025 4.490 127.175 ;
        RECT 0.985 125.220 6.000 127.025 ;
        RECT 0.985 121.925 4.490 125.220 ;
        RECT 0.985 121.115 4.485 121.925 ;
        RECT 0.985 120.965 4.490 121.115 ;
        RECT 0.985 119.160 6.000 120.965 ;
        RECT 0.985 115.865 4.490 119.160 ;
        RECT 0.985 87.265 4.485 115.865 ;
        RECT 296.815 114.965 300.315 220.405 ;
        RECT 295.300 114.355 300.315 114.965 ;
        RECT 296.815 112.405 300.315 114.355 ;
        RECT 295.300 111.810 300.315 112.405 ;
        RECT 296.815 87.265 300.315 111.810 ;
        RECT 0.985 86.795 6.000 87.265 ;
        RECT 295.300 86.795 300.315 87.265 ;
        RECT 0.985 72.515 4.485 86.795 ;
        RECT 296.815 72.515 300.315 86.795 ;
        RECT 0.985 71.835 6.000 72.515 ;
        RECT 295.300 71.835 300.315 72.515 ;
        RECT 0.985 4.485 4.485 71.835 ;
        RECT 95.850 4.485 202.075 6.000 ;
        RECT 296.815 4.485 300.315 71.835 ;
        RECT 0.985 4.480 202.505 4.485 ;
        RECT 204.680 4.480 300.315 4.485 ;
        RECT 0.985 0.985 300.315 4.480 ;
        RECT 87.030 0.980 87.730 0.985 ;
        RECT 90.590 0.980 91.290 0.985 ;
      LAYER Metal2 ;
        RECT 0.985 222.800 300.315 223.940 ;
        RECT 0.995 215.810 2.125 218.240 ;
        RECT 299.120 215.795 300.800 218.225 ;
        RECT 0.995 209.750 2.125 212.180 ;
        RECT 299.120 209.735 300.800 212.165 ;
        RECT 0.995 203.690 2.125 206.120 ;
        RECT 299.120 203.675 300.800 206.105 ;
        RECT 0.995 197.630 2.125 200.060 ;
        RECT 299.120 197.615 300.800 200.045 ;
        RECT 0.995 191.570 2.125 194.000 ;
        RECT 299.120 191.555 300.800 193.985 ;
        RECT 0.995 185.510 2.125 187.940 ;
        RECT 299.120 185.495 300.800 187.925 ;
        RECT 0.995 179.450 2.125 181.880 ;
        RECT 299.120 179.435 300.800 181.865 ;
        RECT 0.995 173.390 2.125 175.820 ;
        RECT 299.120 173.375 300.800 175.805 ;
        RECT 0.995 167.330 2.125 169.760 ;
        RECT 299.120 167.315 300.800 169.745 ;
        RECT 0.995 161.270 2.125 163.700 ;
        RECT 299.120 161.255 300.800 163.685 ;
        RECT 0.995 155.210 2.125 157.640 ;
        RECT 299.120 155.195 300.800 157.625 ;
        RECT 0.995 149.150 2.125 151.580 ;
        RECT 299.120 149.135 300.800 151.565 ;
        RECT 0.995 143.090 2.125 145.520 ;
        RECT 299.120 143.075 300.800 145.505 ;
        RECT 0.995 137.030 2.125 139.460 ;
        RECT 299.120 137.015 300.800 139.445 ;
        RECT 0.995 130.970 2.125 133.400 ;
        RECT 299.120 130.955 300.800 133.385 ;
        RECT 0.995 124.910 2.125 127.340 ;
        RECT 299.120 124.895 300.800 127.325 ;
        RECT 0.995 118.850 2.125 121.280 ;
        RECT 299.120 118.835 300.800 121.265 ;
        RECT 0.995 111.495 2.125 113.925 ;
        RECT 299.185 111.495 300.315 113.925 ;
        RECT 0.995 83.455 2.125 92.695 ;
        RECT 299.185 83.455 300.315 92.695 ;
        RECT 0.995 69.460 2.125 72.760 ;
        RECT 299.185 69.460 300.315 72.760 ;
        RECT 0.995 48.095 2.125 57.145 ;
        RECT 299.185 48.095 300.315 57.145 ;
        RECT 0.995 33.790 2.125 37.960 ;
        RECT 299.185 33.790 300.315 37.960 ;
        RECT 0.995 19.880 2.125 26.220 ;
        RECT 299.185 19.880 300.315 26.220 ;
        RECT 0.995 8.890 2.125 13.060 ;
        RECT 299.185 8.890 300.315 13.060 ;
        RECT 16.245 0.985 19.745 4.485 ;
        RECT 25.040 0.985 25.820 6.000 ;
        RECT 28.600 0.985 29.385 6.000 ;
        RECT 33.045 0.985 36.545 4.485 ;
        RECT 54.045 0.985 57.545 4.485 ;
        RECT 63.850 0.985 64.630 6.000 ;
        RECT 67.410 0.985 68.195 6.000 ;
        RECT 70.845 0.985 74.345 4.485 ;
        RECT 87.000 0.975 87.775 6.000 ;
        RECT 90.555 0.975 91.335 6.000 ;
        RECT 101.350 4.800 102.480 6.000 ;
        RECT 101.520 1.450 102.305 4.800 ;
        RECT 109.630 0.985 113.130 4.485 ;
        RECT 115.575 0.985 119.075 4.485 ;
        RECT 121.905 0.985 125.405 4.485 ;
        RECT 129.495 4.310 130.275 6.000 ;
        RECT 133.055 4.485 133.840 6.000 ;
        RECT 135.865 4.485 136.645 6.000 ;
        RECT 133.055 4.310 136.645 4.485 ;
        RECT 139.425 4.310 140.210 6.000 ;
        RECT 133.095 0.985 136.595 4.310 ;
        RECT 144.315 0.985 147.815 4.485 ;
        RECT 152.715 0.985 156.215 4.485 ;
        RECT 161.115 0.985 164.615 4.485 ;
        RECT 179.315 0.985 182.815 4.485 ;
        RECT 183.670 0.985 187.170 4.485 ;
        RECT 206.100 1.005 206.875 6.000 ;
        RECT 209.655 1.005 210.435 6.000 ;
        RECT 223.760 0.985 227.260 4.485 ;
        RECT 230.315 0.985 231.095 6.000 ;
        RECT 233.875 0.985 234.660 6.000 ;
        RECT 240.560 0.985 244.060 4.485 ;
        RECT 261.560 0.985 265.060 4.485 ;
        RECT 269.465 0.965 270.245 6.000 ;
        RECT 273.025 0.965 273.810 6.000 ;
        RECT 278.360 0.985 281.860 4.485 ;
      LAYER Metal3 ;
        RECT 9.370 222.795 12.870 224.930 ;
        RECT 18.760 222.800 22.260 224.930 ;
        RECT 28.910 222.795 32.410 224.930 ;
        RECT 37.660 222.800 41.160 224.930 ;
        RECT 48.450 222.795 51.950 224.930 ;
        RECT 56.560 222.800 60.060 224.930 ;
        RECT 67.990 222.795 71.490 224.930 ;
        RECT 80.400 222.795 83.900 224.930 ;
        RECT 88.805 222.800 92.305 224.930 ;
        RECT 98.320 222.800 101.820 224.930 ;
        RECT 103.205 222.800 106.705 224.930 ;
        RECT 114.085 222.800 117.585 224.930 ;
        RECT 119.835 222.800 123.335 224.930 ;
        RECT 130.070 222.800 133.570 224.930 ;
        RECT 140.340 222.800 143.840 224.930 ;
        RECT 149.255 222.800 152.755 224.930 ;
        RECT 153.745 222.800 157.245 224.930 ;
        RECT 166.375 222.800 169.875 224.930 ;
        RECT 177.380 222.800 180.880 224.930 ;
        RECT 196.715 222.800 200.215 224.930 ;
        RECT 205.520 222.800 209.020 224.930 ;
        RECT 214.800 222.795 218.300 224.930 ;
        RECT 226.275 222.800 229.775 224.930 ;
        RECT 234.340 222.795 237.840 224.930 ;
        RECT 245.175 222.800 248.675 224.930 ;
        RECT 253.880 222.795 257.380 224.930 ;
        RECT 264.075 222.800 267.575 224.930 ;
        RECT 273.420 222.795 276.920 224.930 ;
        RECT 285.830 222.795 289.330 224.930 ;
        RECT 0.000 217.550 3.555 218.250 ;
        RECT 297.755 218.130 301.300 218.235 ;
        RECT 297.750 217.735 301.300 218.130 ;
        RECT 0.000 216.500 6.000 217.550 ;
        RECT 295.300 216.685 301.300 217.735 ;
        RECT 0.000 215.800 3.555 216.500 ;
        RECT 297.750 215.685 301.300 216.685 ;
        RECT 0.000 211.490 3.555 212.190 ;
        RECT 297.750 211.675 301.300 212.175 ;
        RECT 0.000 210.440 6.000 211.490 ;
        RECT 295.300 210.625 301.300 211.675 ;
        RECT 0.000 209.740 3.555 210.440 ;
        RECT 297.750 209.725 301.300 210.625 ;
        RECT 0.000 205.430 3.555 206.130 ;
        RECT 297.750 205.615 301.300 206.115 ;
        RECT 0.000 204.380 6.000 205.430 ;
        RECT 295.300 204.565 301.300 205.615 ;
        RECT 0.000 203.680 3.555 204.380 ;
        RECT 297.750 203.665 301.300 204.565 ;
        RECT 0.000 199.370 3.555 200.070 ;
        RECT 297.750 199.555 301.300 200.055 ;
        RECT 0.000 198.320 6.000 199.370 ;
        RECT 295.300 198.505 301.300 199.555 ;
        RECT 0.000 197.620 3.555 198.320 ;
        RECT 297.750 197.605 301.300 198.505 ;
        RECT 0.000 193.310 3.555 194.010 ;
        RECT 297.750 193.495 301.300 193.995 ;
        RECT 0.000 192.260 6.000 193.310 ;
        RECT 295.300 192.445 301.300 193.495 ;
        RECT 0.000 191.560 3.555 192.260 ;
        RECT 297.750 191.545 301.300 192.445 ;
        RECT 0.000 187.250 3.555 187.950 ;
        RECT 297.750 187.435 301.300 187.935 ;
        RECT 0.000 186.200 6.000 187.250 ;
        RECT 295.300 186.385 301.300 187.435 ;
        RECT 0.000 185.500 3.555 186.200 ;
        RECT 297.750 185.485 301.300 186.385 ;
        RECT 0.000 181.190 3.555 181.890 ;
        RECT 297.750 181.375 301.300 181.875 ;
        RECT 0.000 180.140 6.000 181.190 ;
        RECT 295.300 180.325 301.300 181.375 ;
        RECT 0.000 179.440 3.555 180.140 ;
        RECT 297.750 179.425 301.300 180.325 ;
        RECT 0.000 175.130 3.555 175.830 ;
        RECT 297.750 175.315 301.300 175.815 ;
        RECT 0.000 174.080 6.000 175.130 ;
        RECT 295.300 174.265 301.300 175.315 ;
        RECT 0.000 173.380 3.555 174.080 ;
        RECT 297.750 173.365 301.300 174.265 ;
        RECT 0.000 169.070 3.555 169.770 ;
        RECT 297.750 169.255 301.300 169.755 ;
        RECT 0.000 168.020 6.000 169.070 ;
        RECT 295.300 168.205 301.300 169.255 ;
        RECT 0.000 167.320 3.555 168.020 ;
        RECT 297.750 167.305 301.300 168.205 ;
        RECT 0.000 163.010 3.555 163.710 ;
        RECT 297.750 163.195 301.300 163.695 ;
        RECT 0.000 161.960 6.000 163.010 ;
        RECT 295.300 162.145 301.300 163.195 ;
        RECT 0.000 161.260 3.555 161.960 ;
        RECT 297.750 161.245 301.300 162.145 ;
        RECT 0.000 156.950 3.555 157.650 ;
        RECT 297.750 157.135 301.300 157.635 ;
        RECT 0.000 155.900 6.000 156.950 ;
        RECT 295.300 156.085 301.300 157.135 ;
        RECT 0.000 155.200 3.555 155.900 ;
        RECT 297.750 155.185 301.300 156.085 ;
        RECT 0.000 150.890 3.555 151.590 ;
        RECT 297.750 151.075 301.300 151.575 ;
        RECT 0.000 149.840 6.000 150.890 ;
        RECT 295.300 150.025 301.300 151.075 ;
        RECT 0.000 149.140 3.555 149.840 ;
        RECT 297.750 149.125 301.300 150.025 ;
        RECT 0.000 144.830 3.555 145.530 ;
        RECT 297.750 145.015 301.300 145.515 ;
        RECT 0.000 143.780 6.000 144.830 ;
        RECT 295.300 143.965 301.300 145.015 ;
        RECT 0.000 143.080 3.555 143.780 ;
        RECT 297.750 143.065 301.300 143.965 ;
        RECT 0.000 138.770 3.555 139.470 ;
        RECT 297.750 138.955 301.300 139.455 ;
        RECT 0.000 137.720 6.000 138.770 ;
        RECT 295.300 137.905 301.300 138.955 ;
        RECT 0.000 137.020 3.555 137.720 ;
        RECT 297.750 137.005 301.300 137.905 ;
        RECT 0.000 132.710 3.555 133.410 ;
        RECT 297.750 132.895 301.300 133.395 ;
        RECT 0.000 131.660 6.000 132.710 ;
        RECT 295.300 131.845 301.300 132.895 ;
        RECT 0.000 130.960 3.555 131.660 ;
        RECT 297.750 130.945 301.300 131.845 ;
        RECT 0.000 126.650 3.555 127.350 ;
        RECT 297.755 127.190 301.300 127.335 ;
        RECT 297.750 126.835 301.300 127.190 ;
        RECT 0.000 125.600 6.000 126.650 ;
        RECT 295.300 125.785 301.300 126.835 ;
        RECT 0.000 124.900 3.555 125.600 ;
        RECT 297.750 124.885 301.300 125.785 ;
        RECT 0.000 120.590 3.555 121.290 ;
        RECT 297.755 121.080 301.300 121.275 ;
        RECT 297.750 120.775 301.300 121.080 ;
        RECT 0.000 119.540 6.000 120.590 ;
        RECT 295.300 119.725 301.300 120.775 ;
        RECT 0.000 118.840 3.555 119.540 ;
        RECT 297.750 118.825 301.300 119.725 ;
        RECT 0.010 114.115 6.000 114.360 ;
        RECT 0.000 113.660 6.000 114.115 ;
        RECT 295.300 113.660 301.300 114.360 ;
        RECT 0.000 113.025 3.555 113.660 ;
        RECT 297.750 113.025 301.300 113.660 ;
        RECT 0.000 111.350 6.000 113.025 ;
        RECT 0.010 111.345 6.000 111.350 ;
        RECT 295.300 111.345 301.300 113.025 ;
        RECT 0.000 93.825 3.545 93.830 ;
        RECT 297.750 93.825 301.300 93.830 ;
        RECT 0.000 86.895 6.000 93.825 ;
        RECT 0.010 86.890 6.000 86.895 ;
        RECT 295.300 86.890 301.300 93.825 ;
        RECT 295.300 86.830 295.500 86.890 ;
        RECT 0.000 72.855 0.700 72.860 ;
        RECT 297.755 72.855 301.300 72.860 ;
        RECT 0.000 71.265 6.000 72.855 ;
        RECT 295.300 71.265 301.300 72.855 ;
        RECT 0.000 69.355 3.555 71.265 ;
        RECT 297.755 70.860 301.300 71.265 ;
        RECT 297.750 69.355 301.300 70.860 ;
        RECT 0.000 47.950 6.000 57.210 ;
        RECT 295.300 47.950 301.300 57.210 ;
        RECT 297.750 38.225 301.300 38.230 ;
        RECT 0.000 33.615 6.000 38.225 ;
        RECT 295.300 33.615 301.300 38.225 ;
        RECT 0.000 23.645 6.000 25.465 ;
        RECT 295.300 23.645 301.300 25.465 ;
        RECT 0.000 23.315 3.565 23.645 ;
        RECT 297.745 23.315 301.300 23.645 ;
        RECT 0.000 21.325 3.555 23.315 ;
        RECT 297.750 21.325 301.300 23.315 ;
        RECT 0.000 19.810 6.000 21.325 ;
        RECT 295.300 19.810 301.300 21.325 ;
        RECT 0.000 13.195 0.700 13.200 ;
        RECT 0.000 11.965 6.000 13.195 ;
        RECT 295.300 11.965 301.300 13.195 ;
        RECT 0.000 9.985 3.545 11.965 ;
        RECT 297.805 9.985 301.300 11.965 ;
        RECT 0.000 8.740 6.000 9.985 ;
        RECT 295.300 8.750 301.300 9.985 ;
        RECT 295.300 8.745 298.065 8.750 ;
        RECT 16.245 0.000 19.745 3.260 ;
        RECT 33.045 0.000 36.545 3.260 ;
        RECT 54.045 0.000 57.545 3.260 ;
        RECT 70.845 0.000 74.345 3.260 ;
        RECT 109.630 0.000 113.130 3.260 ;
        RECT 115.575 0.000 119.075 3.260 ;
        RECT 121.905 0.000 125.405 3.260 ;
        RECT 133.095 0.000 136.595 3.260 ;
        RECT 144.315 0.000 147.815 3.260 ;
        RECT 152.715 0.000 156.215 3.260 ;
        RECT 161.115 0.000 164.615 3.260 ;
        RECT 179.315 0.000 182.815 3.260 ;
        RECT 183.670 0.000 187.170 3.260 ;
        RECT 223.760 0.000 227.260 3.260 ;
        RECT 240.560 0.000 244.060 3.260 ;
        RECT 261.560 0.000 265.060 3.260 ;
        RECT 278.360 0.000 281.860 3.260 ;
    END
  END VSS
  PIN WEN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 288.510 5.985 289.140 5.990 ;
        RECT 288.510 5.955 289.420 5.985 ;
        RECT 288.510 5.695 290.025 5.955 ;
        RECT 288.510 5.685 289.420 5.695 ;
        RECT 288.510 5.650 289.140 5.685 ;
      LAYER Metal2 ;
        RECT 288.430 0.000 289.215 5.995 ;
    END
  END WEN[7]
  PIN WEN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 253.790 5.985 254.350 5.995 ;
        RECT 253.285 5.965 254.350 5.985 ;
        RECT 253.185 5.705 254.355 5.965 ;
        RECT 253.285 5.695 254.350 5.705 ;
        RECT 253.285 5.645 253.915 5.695 ;
      LAYER Metal2 ;
        RECT 253.205 0.000 253.985 6.000 ;
    END
  END WEN[6]
  PIN WEN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 249.780 5.950 250.340 5.980 ;
        RECT 250.710 5.950 251.340 5.985 ;
        RECT 249.775 5.690 251.340 5.950 ;
        RECT 249.780 5.680 250.340 5.690 ;
        RECT 250.710 5.645 251.340 5.690 ;
      LAYER Metal2 ;
        RECT 250.630 0.000 251.410 6.000 ;
    END
  END WEN[5]
  PIN WEN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 214.105 5.950 215.275 5.990 ;
        RECT 214.105 5.690 217.180 5.950 ;
        RECT 216.480 5.600 217.110 5.690 ;
      LAYER Metal2 ;
        RECT 216.400 0.000 217.185 5.955 ;
    END
  END WEN[4]
  PIN WEN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 81.990 5.975 82.620 5.990 ;
        RECT 83.305 5.975 83.865 5.980 ;
        RECT 81.950 5.950 84.110 5.975 ;
        RECT 81.950 5.690 84.470 5.950 ;
        RECT 81.950 5.670 84.110 5.690 ;
        RECT 81.990 5.650 82.620 5.670 ;
      LAYER Metal2 ;
        RECT 81.910 0.000 82.695 6.000 ;
    END
  END WEN[3]
  PIN WEN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 45.915 5.940 46.545 5.990 ;
        RECT 48.235 5.960 48.795 5.990 ;
        RECT 47.630 5.940 48.800 5.960 ;
        RECT 45.915 5.700 48.800 5.940 ;
        RECT 45.915 5.690 48.795 5.700 ;
        RECT 45.915 5.665 48.390 5.690 ;
        RECT 45.915 5.650 46.545 5.665 ;
      LAYER Metal2 ;
        RECT 45.685 5.650 46.545 5.990 ;
        RECT 45.685 0.000 46.470 5.650 ;
    END
  END WEN[2]
  PIN WEN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 44.190 5.980 44.820 5.990 ;
        RECT 44.190 5.950 45.035 5.980 ;
        RECT 44.190 5.690 45.640 5.950 ;
        RECT 44.190 5.680 45.035 5.690 ;
        RECT 44.190 5.665 44.945 5.680 ;
        RECT 44.190 5.650 44.820 5.665 ;
      LAYER Metal2 ;
        RECT 44.110 0.000 44.895 5.995 ;
    END
  END WEN[1]
  PIN WEN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.800 5.650 10.850 6.000 ;
        RECT 10.215 5.645 10.845 5.650 ;
      LAYER Metal2 ;
        RECT 10.215 5.980 10.845 5.985 ;
        RECT 10.085 0.000 10.870 5.980 ;
    END
  END WEN[0]
  OBS
      LAYER Nwell ;
        RECT 6.305 6.000 295.010 218.930 ;
      LAYER Metal1 ;
        RECT 6.000 6.000 295.300 218.930 ;
      LAYER Metal2 ;
        RECT 6.000 6.000 295.300 218.930 ;
      LAYER Metal3 ;
        RECT 6.000 86.350 295.300 218.930 ;
        RECT 6.000 85.600 295.500 86.350 ;
        RECT 6.000 85.125 295.300 85.600 ;
        RECT 6.000 84.370 295.500 85.125 ;
        RECT 6.000 83.900 295.300 84.370 ;
        RECT 6.000 83.145 295.500 83.900 ;
        RECT 6.000 82.675 295.300 83.145 ;
        RECT 6.000 81.920 295.500 82.675 ;
        RECT 6.000 6.000 295.300 81.920 ;
  END
END gf180mcu_ocd_ip_sram__sram256x8m8wm1
END LIBRARY

