magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< psubdiff >>
rect -118 23 111 57
rect -118 -23 -78 23
rect 78 -23 111 23
rect -118 -58 111 -23
<< psubdiffcont >>
rect -78 -23 78 23
<< metal1 >>
rect -118 23 105 51
rect -118 -23 -78 23
rect 78 -23 105 23
rect -118 -51 105 -23
<< end >>
