magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< polysilicon >>
rect -181 211 -126 245
rect -22 211 34 245
rect 140 211 196 245
rect 300 211 356 245
rect 462 211 518 245
rect 622 211 678 245
rect 784 211 840 245
rect -181 -34 -126 0
rect -22 -34 34 0
rect 140 -34 196 0
rect 300 -34 356 0
rect 462 -34 518 0
rect 622 -34 678 0
rect 784 -34 840 0
use nmos_5p04310591302026_3v512x8m81  nmos_5p04310591302026_3v512x8m81_0
timestamp 1763765945
transform 1 0 -14 0 1 0
box -256 -44 942 255
<< end >>
