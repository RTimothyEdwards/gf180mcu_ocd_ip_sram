magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< psubdiff >>
rect -55 194 56 228
rect -55 -194 -23 194
rect 23 -194 56 194
rect -55 -228 56 -194
<< psubdiffcont >>
rect -23 -194 23 194
<< metal1 >>
rect -49 194 49 222
rect -49 -194 -23 194
rect 23 -194 49 194
rect -49 -222 49 -194
<< end >>
