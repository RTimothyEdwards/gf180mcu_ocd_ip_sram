magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal1 >>
rect -119 322 119 351
rect -119 -322 -92 322
rect 92 -322 119 322
rect -119 -351 119 -322
<< via1 >>
rect -92 -322 92 322
<< metal2 >>
rect -119 322 119 351
rect -119 -322 -92 322
rect 92 -322 119 322
rect -119 -351 119 -322
<< end >>
