magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal1 >>
rect -44 102 45 123
rect -44 -102 -26 102
rect 26 -102 45 102
rect -44 -122 45 -102
<< via1 >>
rect -26 -102 26 102
<< metal2 >>
rect -45 102 45 123
rect -45 -102 -26 102
rect 26 -102 45 102
rect -45 -123 45 -102
<< end >>
