magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< psubdiff >>
rect -1383 130 1383 172
rect -1383 -130 -1344 130
rect 1344 -130 1383 130
rect -1383 -171 1383 -130
<< psubdiffcont >>
rect -1344 -130 1344 130
<< metal1 >>
rect -1378 130 1377 165
rect -1378 -130 -1344 130
rect 1344 -130 1377 130
rect -1378 -165 1377 -130
<< end >>
