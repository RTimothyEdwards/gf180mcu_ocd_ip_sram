magic
tech gf180mcuD
magscale 1 10
timestamp 1763486358
<< nwell >>
rect 3794 18861 3871 19309
rect 4879 18886 5119 19213
rect 8943 18861 9012 19309
rect 9991 18886 10273 19213
rect 17413 18886 18305 19293
rect 2429 14978 2450 16568
rect 6305 15569 6363 17303
rect 7591 14978 7617 16568
rect 16172 15253 16226 16836
rect 3842 12864 6164 13696
rect 9007 12864 11329 13696
rect 4106 12863 4203 12864
rect 5286 12863 5386 12864
rect 9274 12863 9367 12864
rect 10456 12863 10547 12864
rect 17262 6999 17293 7020
rect 18106 6999 18193 7020
rect 18983 6999 19055 7020
rect 14494 5649 15036 6010
rect 16382 5953 19055 6999
rect 14517 4696 14632 4729
rect 17262 4106 17293 5953
rect 18106 3677 18193 5953
rect 18983 3771 19055 5953
rect 5846 504 6015 912
<< metal1 >>
rect 282 808 375 20325
rect 1143 20257 1270 20304
rect 4808 12337 4899 12478
rect 535 12243 4899 12337
rect 535 7506 625 12243
rect 6001 12178 6092 12469
rect 704 12084 6092 12178
rect 704 7770 795 12084
rect 9952 12019 10042 12457
rect 873 11926 10042 12019
rect 11136 12073 11226 12511
rect 17292 12232 17383 12523
rect 18476 12391 18566 12532
rect 19649 12456 20202 12549
rect 18476 12297 20033 12391
rect 17292 12139 19864 12232
rect 11136 11980 19695 12073
rect 873 7975 963 11926
rect 873 7886 1290 7975
rect 704 7661 1121 7770
rect 535 7399 952 7506
rect 861 564 952 7399
rect 1031 564 1121 7661
rect 1199 564 1290 7886
rect 14693 6741 14743 6870
rect 15017 6741 15068 6875
rect 15336 6741 15386 6861
rect 14693 6691 15386 6741
rect 14710 6690 15369 6691
rect 15701 1162 15748 1164
rect 14532 1113 15748 1162
rect 9200 285 10308 333
rect 15701 307 15748 1113
rect 19604 421 19695 11980
rect 19773 421 19864 12139
rect 19943 421 20033 12297
rect 20111 421 20202 12456
rect 20664 808 20757 20325
rect 282 -88 6454 231
rect 9200 -1052 9248 285
rect 19488 -88 20590 231
<< metal2 >>
rect 451 967 1043 21087
rect 12009 20205 12100 20298
rect 12255 20205 12345 20298
rect 13153 20205 13244 20298
rect 13402 20205 13492 20298
rect 14298 20205 14389 20298
rect 14538 20205 14628 20298
rect 15439 20205 15529 20298
rect 15691 20205 15781 20298
rect 1635 20046 1725 20140
rect 1883 20046 1974 20140
rect 2887 20046 2978 20140
rect 3141 20046 3231 20140
rect 6799 20046 6890 20140
rect 7049 20046 7139 20140
rect 8052 20046 8143 20140
rect 8306 20046 8397 20140
rect 6274 1224 6364 1376
rect 5693 1130 6364 1224
rect 11423 1155 11480 1157
rect 282 -998 375 809
rect 451 -88 760 967
rect 861 -998 952 809
rect 1031 -998 1121 809
rect 1199 -998 1290 809
rect 2359 -998 2452 1062
rect 3542 -998 3636 1062
rect 4727 -998 4821 1062
rect 5693 -692 5783 1130
rect 11353 1116 11480 1155
rect 6216 116 6454 1024
rect 11423 -956 11480 1116
rect 15128 -100 15375 2419
rect 19972 967 20588 21087
rect 15998 -998 16092 432
rect 19604 -998 19695 819
rect 19773 -998 19864 819
rect 19943 -998 20033 819
rect 20111 -998 20202 819
rect 20279 -88 20588 967
rect 20664 -880 20757 809
<< metal3 >>
rect 451 20451 20588 21087
rect 282 20080 20757 20325
rect 19677 10387 19767 10480
rect 19677 10149 19767 10242
rect 19677 9911 19767 10004
rect 19677 9673 19767 9766
rect 19677 9435 19767 9528
rect 19677 9197 19767 9290
rect 19677 8958 19767 9052
rect 19677 8720 19767 8814
rect 9743 4890 9967 5501
use gen_512x8_512x8m81  gen_512x8_512x8m81_0
timestamp 1763486358
transform 1 0 9916 0 1 499
box -12453 -1374 12336 11499
use M1_NACTIVE4310591302047_512x8m81  M1_NACTIVE4310591302047_512x8m81_0
timestamp 1763476864
transform 0 -1 18221 1 0 19080
box -62 -36 62 36
use M1_NACTIVE4310591302047_512x8m81  M1_NACTIVE4310591302047_512x8m81_1
timestamp 1763476864
transform 0 -1 17500 1 0 19119
box -62 -36 62 36
use M1_PACTIVE4310591302048_512x8m81  M1_PACTIVE4310591302048_512x8m81_0
timestamp 1763476864
transform 1 0 2440 0 1 20281
box -1113 -36 1153 36
use M1_PACTIVE4310591302048_512x8m81  M1_PACTIVE4310591302048_512x8m81_1
timestamp 1763476864
transform 1 0 7592 0 1 20281
box -1113 -36 1153 36
use M1_PACTIVE4310591302049_512x8m81  M1_PACTIVE4310591302049_512x8m81_0
timestamp 1763476864
transform 1 0 16713 0 1 19868
box -457 -36 457 36
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1763476864
transform -1 0 20710 0 1 20202
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_1
timestamp 1763476864
transform -1 0 20710 0 1 687
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_2
timestamp 1763476864
transform 1 0 329 0 1 20202
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_3
timestamp 1763476864
transform 1 0 329 0 1 687
box -43 -122 43 122
use M2_M1$$199746604_512x8m81  M2_M1$$199746604_512x8m81_0
timestamp 1763476864
transform 1 0 605 0 1 71
box -119 -123 119 123
use M2_M1$$199746604_512x8m81  M2_M1$$199746604_512x8m81_1
timestamp 1763476864
transform 1 0 20433 0 1 71
box -119 -123 119 123
use M2_M1$$199746604_512x8m81  M2_M1$$199746604_512x8m81_2
timestamp 1763476864
transform 1 0 6335 0 1 -3
box -119 -123 119 123
use M2_M1$$201262124_512x8m81  M2_M1$$201262124_512x8m81_0
timestamp 1763476864
transform 1 0 6335 0 1 184
box -119 -46 119 46
use M2_M1$$202405932_512x8m81  M2_M1$$202405932_512x8m81_0
timestamp 1763476864
transform 1 0 20157 0 1 620
box -44 -198 44 198
use M2_M1$$202405932_512x8m81  M2_M1$$202405932_512x8m81_1
timestamp 1763476864
transform 1 0 19988 0 1 620
box -44 -198 44 198
use M2_M1$$202405932_512x8m81  M2_M1$$202405932_512x8m81_2
timestamp 1763476864
transform 1 0 19819 0 1 620
box -44 -198 44 198
use M2_M1$$202405932_512x8m81  M2_M1$$202405932_512x8m81_3
timestamp 1763476864
transform 1 0 19649 0 1 620
box -44 -198 44 198
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_0
timestamp 1763476864
transform 1 0 1245 0 1 687
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_1
timestamp 1763476864
transform 1 0 1075 0 1 687
box -45 -122 45 123
use M2_M1$$202406956_512x8m81  M2_M1$$202406956_512x8m81_2
timestamp 1763476864
transform 1 0 907 0 1 687
box -45 -122 45 123
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_0
timestamp 1763476864
transform -1 0 20710 0 1 20202
box -44 -123 44 123
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_1
timestamp 1763476864
transform 1 0 329 0 1 20202
box -44 -123 44 123
use M3_M2$$201255980_512x8m81  M3_M2$$201255980_512x8m81_0
timestamp 1763476864
transform -1 0 20640 0 1 -672
box -119 -46 119 46
use M3_M2$$201255980_512x8m81  M3_M2$$201255980_512x8m81_1
timestamp 1763476864
transform 1 0 399 0 1 -672
box -119 -46 119 46
use M3_M2$$201255980_512x8m81  M3_M2$$201255980_512x8m81_2
timestamp 1763476864
transform 1 0 5738 0 1 -672
box -119 -46 119 46
use M3_M2$$201401388_512x8m81  M3_M2$$201401388_512x8m81_0
timestamp 1763476864
transform 1 0 20280 0 1 20769
box -266 -275 266 275
use M3_M2$$201401388_512x8m81  M3_M2$$201401388_512x8m81_1
timestamp 1763476864
transform 1 0 759 0 1 20769
box -266 -275 266 275
use M3_M2$$201401388_512x8m81  M3_M2$$201401388_512x8m81_2
timestamp 1763476864
transform 1 0 20280 0 1 6782
box -266 -275 266 275
use M3_M24310591302050_512x8m81  M3_M24310591302050_512x8m81_0
timestamp 1763476864
transform 1 0 15254 0 1 56
box -99 -99 99 99
use M3_M24310591302050_512x8m81  M3_M24310591302050_512x8m81_1
timestamp 1763476864
transform 1 0 15254 0 1 672
box -99 -99 99 99
use prexdec_top_512x8m81  prexdec_top_512x8m81_0
timestamp 1763476864
transform 1 0 949 0 1 12306
box 21 -1 19120 8780
use ypredec1_512x8m81  ypredec1_512x8m81_0
timestamp 1763476864
transform 1 0 1092 0 1 392
box 125 53 18674 11572
<< labels >>
flabel metal3 s 5796 -700 5796 -700 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 5796 -246 5796 -246 0 FreeSans 313 0 0 0 VDD
port 2 nsew
rlabel metal3 s 19722 10434 19722 10434 4 RYS[7]
port 3 nsew
rlabel metal3 s 19722 10195 19722 10195 4 RYS[6]
port 4 nsew
rlabel metal3 s 19722 9957 19722 9957 4 RYS[5]
port 5 nsew
rlabel metal3 s 19722 9719 19722 9719 4 RYS[4]
port 6 nsew
rlabel metal3 s 19722 9481 19722 9481 4 RYS[3]
port 7 nsew
rlabel metal3 s 19722 9243 19722 9243 4 RYS[2]
port 8 nsew
rlabel metal3 s 19722 9005 19722 9005 4 RYS[1]
port 9 nsew
rlabel metal3 s 19722 8767 19722 8767 4 RYS[0]
port 10 nsew
rlabel metal3 s 1263 8767 1263 8767 4 LYS[0]
port 11 nsew
rlabel metal3 s 1263 9005 1263 9005 4 LYS[1]
port 12 nsew
rlabel metal3 s 1263 9243 1263 9243 4 LYS[2]
port 13 nsew
rlabel metal3 s 1263 9481 1263 9481 4 LYS[3]
port 14 nsew
rlabel metal3 s 1263 10195 1263 10195 4 LYS[6]
port 15 nsew
rlabel metal3 s 1263 9957 1263 9957 4 LYS[5]
port 16 nsew
rlabel metal3 s 1263 9719 1263 9719 4 LYS[4]
port 17 nsew
rlabel metal3 s 18802 20769 18802 20769 4 men
port 18 nsew
rlabel metal3 s 1263 10434 1263 10434 4 LYS[7]
port 19 nsew
rlabel metal3 s 19569 3513 19569 3513 4 tblhl
port 20 nsew
flabel metal3 s 4365 6314 4365 6314 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 4365 12712 4365 12712 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 4365 2449 4365 2449 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 4365 976 4365 976 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 5796 741 5796 741 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 4365 13286 4365 13286 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 4365 16804 4365 16804 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 4365 1713 4365 1713 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 4365 19672 4365 19672 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 4365 18246 4365 18246 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 4365 4577 4365 4577 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 4365 11179 4365 11179 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 4365 18978 4365 18978 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 4365 14201 4365 14201 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal2 s 11449 -938 11449 -938 0 FreeSans 700 0 0 0 IGWEN
port 21 nsew
rlabel metal2 s 6808 20123 6808 20123 4 xb[3]
port 22 nsew
rlabel metal2 s 7114 20128 7114 20128 4 xb[2]
port 23 nsew
rlabel metal2 s 8376 20111 8376 20111 4 xb[0]
port 24 nsew
rlabel metal2 s 12054 20251 12054 20251 4 xa[7]
port 25 nsew
rlabel metal2 s 12300 20251 12300 20251 4 xa[6]
port 26 nsew
rlabel metal2 s 13198 20251 13198 20251 4 xa[5]
port 27 nsew
rlabel metal2 s 13447 20251 13447 20251 4 xa[4]
port 28 nsew
rlabel metal2 s 14343 20251 14343 20251 4 xa[3]
port 29 nsew
rlabel metal2 s 14583 20251 14583 20251 4 xa[2]
port 30 nsew
rlabel metal2 s 4774 -952 4774 -952 4 A[0]
port 31 nsew
rlabel metal2 s 16046 -952 16046 -952 4 CEN
port 32 nsew
rlabel metal2 s 8068 20098 8068 20098 4 xb[1]
port 33 nsew
rlabel metal2 s 7094 20093 7094 20093 4 xb[2]
port 23 nsew
rlabel metal2 s 8351 20090 8351 20090 4 xb[0]
port 24 nsew
rlabel metal2 s 1680 20093 1680 20093 4 xc[3]
port 34 nsew
rlabel metal2 s 2933 20090 2933 20090 4 xc[1]
port 35 nsew
rlabel metal2 s 1929 20093 1929 20093 4 xc[2]
port 36 nsew
rlabel metal2 s 3186 20090 3186 20090 4 xc[0]
port 37 nsew
rlabel metal2 s 15736 20251 15736 20251 4 xa[0]
port 38 nsew
rlabel metal2 s 15484 20251 15484 20251 4 xa[1]
port 39 nsew
rlabel metal2 s 907 -952 907 -952 4 A[9]
port 40 nsew
rlabel metal2 s 1245 -952 1245 -952 4 A[7]
port 41 nsew
rlabel metal2 s 329 -952 329 -952 4 CLK
port 42 nsew
rlabel metal2 s 8098 20090 8098 20090 4 xb[1]
port 33 nsew
rlabel metal2 s 6845 20093 6845 20093 4 xb[3]
port 22 nsew
rlabel metal2 s 2405 -952 2405 -952 4 A[2]
port 43 nsew
rlabel metal2 s 3589 -952 3589 -952 4 A[1]
port 44 nsew
rlabel metal2 s 19649 -952 19649 -952 4 A[6]
port 45 nsew
rlabel metal2 s 20157 -952 20157 -952 4 A[3]
port 46 nsew
rlabel metal2 s 19988 -952 19988 -952 4 A[4]
port 47 nsew
rlabel metal2 s 19819 -952 19819 -952 4 A[5]
port 48 nsew
rlabel metal2 s 1075 -952 1075 -952 4 A[8]
port 49 nsew
flabel metal1 s 15717 737 15717 737 0 FreeSans 700 0 0 0 GWE
port 50 nsew
flabel metal1 s 9219 -938 9219 -938 0 FreeSans 700 0 0 0 GWEN
port 51 nsew
<< properties >>
string path 81.095 8.115 81.735 8.115 81.735 -9.165 
<< end >>
