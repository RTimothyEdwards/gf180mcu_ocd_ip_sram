magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect -133 398 265 417
rect -133 394 185 398
rect -133 -57 -53 394
rect -51 -53 185 394
rect 187 -53 265 398
rect -51 -57 265 -53
rect -133 -66 265 -57
<< polysilicon >>
rect -42 351 13 385
rect 118 351 173 385
rect -42 -34 13 0
rect 118 -34 173 0
use pmos_5p04310591302073_512x8m81  pmos_5p04310591302073_512x8m81_0
timestamp 1763476864
transform 1 0 -14 0 1 0
box -202 -86 362 437
<< end >>
