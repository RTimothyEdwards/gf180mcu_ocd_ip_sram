magic
tech gf180mcuD
magscale 1 10
timestamp 1765833244
<< nwell >>
rect -133 -57 240 456
rect 241 -57 369 456
rect -133 -66 369 -57
<< polysilicon >>
rect -70 423 -15 457
rect 90 423 146 457
rect 251 423 307 457
rect -70 -34 -15 0
rect 90 -34 146 0
rect 251 -34 307 0
use pmos_5p04310591302025_3v256x8m81  pmos_5p04310591302025_3v256x8m81_0
timestamp 1765833244
transform 1 0 -14 0 1 0
box -230 -86 495 509
<< end >>
