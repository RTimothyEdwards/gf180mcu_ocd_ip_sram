magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< metal1 >>
rect -108 26 108 33
rect -108 -26 -89 26
rect 89 -26 108 26
rect -108 -34 108 -26
<< via1 >>
rect -89 -26 89 26
<< metal2 >>
rect -95 26 95 46
rect -95 -26 -89 26
rect 89 -26 95 26
rect -95 -46 95 -26
<< end >>
