magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< nmos >>
rect 0 0 56 657
<< ndiff >>
rect -88 644 0 657
rect -88 13 -75 644
rect -29 13 0 644
rect -88 0 0 13
rect 56 644 144 657
rect 56 13 85 644
rect 131 13 144 644
rect 56 0 144 13
<< ndiffc >>
rect -75 13 -29 644
rect 85 13 131 644
<< polysilicon >>
rect 0 657 56 701
rect 0 -44 56 0
<< metal1 >>
rect -75 644 -29 657
rect -75 0 -29 13
rect 85 644 131 657
rect 85 0 131 13
<< labels >>
flabel ndiffc -40 328 -40 328 0 FreeSans 93 0 0 0 S
flabel ndiffc 96 328 96 328 0 FreeSans 93 0 0 0 D
<< end >>
