magic
tech gf180mcuD
magscale 1 10
timestamp 1764700137
<< metal2 >>
rect -35 128 35 135
rect -35 -128 -28 128
rect 28 -128 35 128
rect -35 -135 35 -128
<< via2 >>
rect -28 -128 28 128
<< metal3 >>
rect -35 128 35 135
rect -35 -128 -28 128
rect 28 -128 35 128
rect -35 -135 35 -128
<< end >>
