magic
tech gf180mcuD
magscale 1 10
timestamp 1765924161
<< nwell >>
rect -161 5039 54 8484
rect -121 2318 3694 2520
rect -121 1751 3715 2318
rect -121 1473 739 1751
rect 902 1503 3715 1751
rect 902 1473 3694 1503
rect -121 1104 3694 1473
<< metal1 >>
rect -16 6908 3476 6960
<< metal2 >>
rect 774 1499 845 1710
rect 1689 1495 1750 1707
rect 2591 1495 2652 1699
<< metal3 >>
rect -575 5420 4956 5618
use M1_NACTIVE4310591302028_3v512x8m81  M1_NACTIVE4310591302028_3v512x8m81_0
timestamp 1764623439
transform 1 0 426 0 1 5519
box -122 -181 122 181
use M1_NACTIVE4310591302028_3v512x8m81  M1_NACTIVE4310591302028_3v512x8m81_1
timestamp 1764623439
transform 1 0 1332 0 1 5519
box -122 -181 122 181
use M1_NACTIVE4310591302028_3v512x8m81  M1_NACTIVE4310591302028_3v512x8m81_2
timestamp 1764623439
transform 1 0 2236 0 1 5519
box -122 -181 122 181
use M1_NACTIVE4310591302028_3v512x8m81  M1_NACTIVE4310591302028_3v512x8m81_3
timestamp 1764623439
transform 1 0 3140 0 1 5519
box -122 -181 122 181
use M2_M14310591302018_3v512x8m81  M2_M14310591302018_3v512x8m81_0
timestamp 1764525316
transform 1 0 426 0 1 5519
box -34 -99 34 99
use M2_M14310591302018_3v512x8m81  M2_M14310591302018_3v512x8m81_1
timestamp 1764525316
transform 1 0 1332 0 1 5519
box -34 -99 34 99
use M2_M14310591302018_3v512x8m81  M2_M14310591302018_3v512x8m81_2
timestamp 1764525316
transform 1 0 2236 0 1 5519
box -34 -99 34 99
use M2_M14310591302018_3v512x8m81  M2_M14310591302018_3v512x8m81_3
timestamp 1764525316
transform 1 0 3140 0 1 5519
box -34 -99 34 99
use M2_M14310591302020_3v512x8m81  M2_M14310591302020_3v512x8m81_0
timestamp 1764525316
transform 1 0 809 0 1 1648
box -35 -56 35 55
use M2_M14310591302020_3v512x8m81  M2_M14310591302020_3v512x8m81_2
timestamp 1764525316
transform 1 0 1719 0 1 1648
box -35 -56 35 55
use M2_M14310591302020_3v512x8m81  M2_M14310591302020_3v512x8m81_4
timestamp 1764525316
transform 1 0 2621 0 1 1648
box -35 -56 35 55
use M3_M2431059130201_3v512x8m81  M3_M2431059130201_3v512x8m81_0
timestamp 1764525316
transform 1 0 809 0 1 1581
box -35 -63 35 63
use M3_M2431059130201_3v512x8m81  M3_M2431059130201_3v512x8m81_1
timestamp 1764525316
transform 1 0 1719 0 1 1581
box -35 -63 35 63
use M3_M2431059130201_3v512x8m81  M3_M2431059130201_3v512x8m81_3
timestamp 1764525316
transform 1 0 2621 0 1 1581
box -35 -63 35 63
use M3_M24310591302029_3v512x8m81  M3_M24310591302029_3v512x8m81_0
timestamp 1764525316
transform 1 0 426 0 1 5519
box -35 -99 35 99
use M3_M24310591302029_3v512x8m81  M3_M24310591302029_3v512x8m81_1
timestamp 1764525316
transform 1 0 1332 0 1 5519
box -35 -99 35 99
use M3_M24310591302029_3v512x8m81  M3_M24310591302029_3v512x8m81_2
timestamp 1764525316
transform 1 0 2236 0 1 5519
box -35 -99 35 99
use M3_M24310591302029_3v512x8m81  M3_M24310591302029_3v512x8m81_3
timestamp 1764525316
transform 1 0 3140 0 1 5519
box -35 -99 35 99
use ypass_gate_3v512x8m81  ypass_gate_3v512x8m81_1
timestamp 1765924077
transform -1 0 3190 0 1 -3377
box -130 4011 633 11861
use ypass_gate_3v512x8m81  ypass_gate_3v512x8m81_2
timestamp 1765924077
transform -1 0 2288 0 1 -3377
box -130 4011 633 11861
use ypass_gate_3v512x8m81  ypass_gate_3v512x8m81_3
timestamp 1765924077
transform -1 0 1386 0 1 -3377
box -130 4011 633 11861
use ypass_gate_3v512x8m81  ypass_gate_3v512x8m81_4
timestamp 1765924077
transform 1 0 2180 0 1 -3377
box -130 4011 633 11861
use ypass_gate_3v512x8m81  ypass_gate_3v512x8m81_5
timestamp 1765924077
transform 1 0 1278 0 1 -3377
box -130 4011 633 11861
use ypass_gate_3v512x8m81  ypass_gate_3v512x8m81_6
timestamp 1765924077
transform 1 0 376 0 1 -3377
box -130 4011 633 11861
use ypass_gate_3v512x8m81  ypass_gate_3v512x8m81_7
timestamp 1765924077
transform -1 0 484 0 1 -3377
box -130 4011 633 11861
use ypass_gate_a_3v512x8m81  ypass_gate_a_3v512x8m81_0
timestamp 1765924161
transform 1 0 3090 0 1 -3377
box -130 4017 627 11860
<< end >>
