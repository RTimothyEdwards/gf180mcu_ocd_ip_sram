magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< nwell >>
rect 341 1390 1141 1714
rect 2 772 1140 1390
<< psubdiff >>
rect 77 672 170 706
rect 77 512 100 672
rect 146 512 170 672
rect 77 477 170 512
<< nsubdiff >>
rect 77 1267 170 1292
rect 77 1036 100 1267
rect 146 1036 170 1267
rect 77 910 170 1036
<< psubdiffcont >>
rect 100 512 146 672
<< nsubdiffcont >>
rect 100 1036 146 1267
<< polysilicon >>
rect 527 1637 583 1783
rect 886 1768 942 1784
rect 886 1722 1166 1768
rect 527 1439 583 1488
rect 262 1397 583 1439
rect 887 1415 941 1484
rect 887 1360 963 1415
rect 1107 1233 1166 1722
rect 886 1185 1166 1233
rect 886 1177 942 1185
rect 372 737 716 833
rect 372 625 428 737
rect 532 625 588 737
rect 886 720 1110 762
rect 886 665 942 720
<< metal1 >>
rect 442 1969 1030 2033
rect 442 1519 523 1969
rect 599 1450 680 1615
rect 251 1426 336 1427
rect 251 1362 523 1426
rect 598 1421 680 1450
rect 83 1267 366 1305
rect 83 1036 100 1267
rect 146 1036 366 1267
rect 83 882 366 1036
rect 82 672 176 705
rect 82 512 100 672
rect 146 655 176 672
rect 146 512 366 655
rect 82 472 366 512
rect 442 467 523 1362
rect 802 827 883 1917
rect 959 1523 1030 1969
rect 1098 1681 1179 1765
rect 938 1348 1164 1431
rect 609 744 883 827
rect 801 714 883 744
rect 802 464 883 714
rect 938 601 1015 1143
rect 1094 726 1150 1348
rect 938 517 1032 601
rect 938 464 1015 517
<< metal3 >>
rect 0 1382 1184 1860
rect 0 936 1184 1298
rect -63 409 1184 861
use M1_POLY2_155_512x8m81  M1_POLY2_155_512x8m81_0
timestamp 1763765945
transform 1 0 648 0 1 786
box -67 -48 67 47
use M1_POLY2_155_512x8m81  M1_POLY2_155_512x8m81_1
timestamp 1763765945
transform 1 0 1130 0 1 768
box -67 -48 67 47
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_0
timestamp 1763765945
transform 1 0 1136 0 1 1707
box -36 -80 36 78
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1763765945
transform 1 0 977 0 1 1390
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1763765945
transform 1 0 291 0 1 1407
box -36 -36 36 36
use M1_PSUB$$45110316_512x8m81  M1_PSUB$$45110316_512x8m81_0
timestamp 1763765945
transform 1 0 214 0 1 1896
box -110 -58 111 57
use M2_M1$$43379756_153_512x8m81  M2_M1$$43379756_153_512x8m81_0
timestamp 1763765945
transform 1 0 639 0 1 1148
box -44 -275 44 275
use M2_M1$$43380780_152_512x8m81  M2_M1$$43380780_152_512x8m81_0
timestamp 1763765945
transform 1 0 127 0 1 1119
box -44 -198 45 198
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_0
timestamp 1763765945
transform 1 0 1139 0 1 1696
box -44 -123 44 122
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_1
timestamp 1763765945
transform 1 0 1138 0 1 1309
box -44 -123 44 122
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_2
timestamp 1763765945
transform 1 0 994 0 1 593
box -44 -123 44 122
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_3
timestamp 1763765945
transform 1 0 124 0 1 581
box -44 -123 44 122
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_4
timestamp 1763765945
transform 1 0 639 0 1 1787
box -44 -123 44 122
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_5
timestamp 1763765945
transform 1 0 123 0 1 1787
box -44 -123 44 122
use M2_M1_154_512x8m81  M2_M1_154_512x8m81_6
timestamp 1763765945
transform 1 0 639 0 1 576
box -44 -123 44 122
use M3_M2$$43368492_151_512x8m81  M3_M2$$43368492_151_512x8m81_0
timestamp 1763765945
transform 1 0 639 0 1 581
box -45 -123 45 123
use M3_M2$$43368492_151_512x8m81  M3_M2$$43368492_151_512x8m81_1
timestamp 1763765945
transform 1 0 124 0 1 581
box -45 -123 45 123
use M3_M2$$47108140_149_512x8m81  M3_M2$$47108140_149_512x8m81_0
timestamp 1763765945
transform 1 0 127 0 1 1109
box -45 -178 45 198
use M3_M2$$47108140_149_512x8m81  M3_M2$$47108140_149_512x8m81_1
timestamp 1763765945
transform 1 0 123 0 1 1657
box -45 -178 45 198
use M3_M2$$47108140_149_512x8m81  M3_M2$$47108140_149_512x8m81_2
timestamp 1763765945
transform 1 0 639 0 1 1657
box -45 -178 45 198
use M3_M2$$47333420_150_512x8m81  M3_M2$$47333420_150_512x8m81_0
timestamp 1763765945
transform 1 0 639 0 1 1036
box -45 -105 45 275
use nmos_1p2$$47329324_512x8m81  nmos_1p2$$47329324_512x8m81_0
timestamp 1763765945
transform 1 0 414 0 1 476
box -130 -44 262 213
use nmos_1p2_157_512x8m81  nmos_1p2_157_512x8m81_0
timestamp 1763765945
transform 1 0 900 0 1 472
box -102 -44 130 255
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_0
timestamp 1763765945
transform 1 0 527 0 -1 1915
box -88 -44 144 133
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_1
timestamp 1763765945
transform 1 0 886 0 -1 1915
box -88 -44 144 133
use pmos_1p2$$47331372_512x8m81  pmos_1p2$$47331372_512x8m81_0
timestamp 1763765945
transform 1 0 414 0 1 877
box -216 -86 348 509
use pmos_1p2_160_512x8m81  pmos_1p2_160_512x8m81_0
timestamp 1763765945
transform 1 0 900 0 1 925
box -188 -86 216 297
use pmos_1p2_161_512x8m81  pmos_1p2_161_512x8m81_0
timestamp 1763765945
transform 1 0 900 0 -1 1615
box -188 -86 216 175
use pmos_1p2_161_512x8m81  pmos_1p2_161_512x8m81_1
timestamp 1763765945
transform 1 0 541 0 -1 1615
box -188 -86 216 175
<< labels >>
rlabel metal1 s 1138 1723 1138 1723 4 enb
port 3 nsew
rlabel metal1 s 1142 1442 1142 1442 4 en
port 4 nsew
rlabel metal1 s 991 559 991 559 4 a
port 6 nsew
rlabel metal1 s 483 499 483 499 4 ab
port 5 nsew
rlabel metal3 s 92 673 92 673 4 vss
port 1 nsew
rlabel metal3 s 109 1156 109 1156 4 vdd
port 2 nsew
rlabel metal3 s 141 1597 141 1597 4 vss
port 1 nsew
<< end >>
