magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
use nmos_5p04310591302016_256x8m81  nmos_5p04310591302016_256x8m81_0
timestamp 1763564386
transform 1 0 -14 0 1 0
box -287 -45 1074 363
<< end >>
