magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nwell >>
rect -178 -66 162 277
rect 163 -57 501 277
rect 502 -57 635 277
rect 163 -66 578 -57
<< polysilicon >>
rect -126 211 -71 245
rect 34 211 89 245
rect 195 211 251 245
rect 355 211 410 245
rect 516 211 572 245
rect -126 -34 -71 0
rect 34 -34 89 0
rect 195 -34 251 0
rect 355 -34 410 0
rect 516 -34 572 0
use pmos_5p04310591302024_3v256x8m81  pmos_5p04310591302024_3v256x8m81_0
timestamp 1763766357
transform 1 0 -14 0 1 0
box -286 -86 760 297
<< end >>
