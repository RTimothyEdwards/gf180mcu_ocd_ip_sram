magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal1 >>
rect -119 703 119 732
rect -119 -703 -92 703
rect 92 -703 119 703
rect -119 -732 119 -703
<< via1 >>
rect -92 -703 92 703
<< metal2 >>
rect -119 703 119 732
rect -119 -703 -92 703
rect 92 -703 119 703
rect -119 -732 119 -703
<< end >>
