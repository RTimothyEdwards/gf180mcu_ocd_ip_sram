magic
tech gf180mcuD
magscale 1 10
timestamp 1765484102
<< nwell >>
rect 4608 77715 6692 78362
rect 9694 78170 10581 78373
rect 9694 78116 10808 78170
rect 7130 77721 7550 77772
rect 9695 77726 10808 78116
rect 4608 77680 6273 77715
rect 11564 77693 14760 78342
<< nsubdiff >>
rect 1486 77791 1594 77953
rect 17843 77805 17952 77953
rect 17842 77664 18051 77805
rect 17842 77578 18034 77664
<< polysilicon >>
rect 4589 78040 5251 78096
rect 4589 77964 4661 78040
rect 4485 77936 4661 77964
rect 7730 77956 7969 77964
rect 4485 77908 5251 77936
rect 7730 77908 8050 77956
rect 4592 77880 5251 77908
rect 7879 77900 8050 77908
rect 8358 77900 8451 77956
rect 9564 77921 9637 78219
rect 10754 77956 10826 78258
rect 12782 78040 13445 78096
rect 10713 77900 10826 77956
rect 10908 77901 11108 77956
rect 10908 77900 11028 77901
rect 11423 77900 11928 77957
rect 14707 77956 14779 78097
rect 12782 77880 13445 77936
rect 14707 77900 15356 77956
rect 14707 77880 14779 77900
<< metal1 >>
rect 1486 77851 2811 78246
rect 3026 78026 4435 78297
rect 4537 77946 5359 78030
rect 4537 77903 4618 77946
rect 1404 77791 2811 77851
rect 4368 77819 4618 77903
rect 6521 77903 6602 78119
rect 7969 78004 8339 78283
rect 9471 78189 9828 78283
rect 8404 78005 8919 78053
rect 9456 78005 10160 78053
rect 10687 77985 10961 78031
rect 11028 77981 11398 78283
rect 11659 78144 14659 78228
rect 11659 78015 12581 78144
rect 12788 77903 12849 78072
rect 14628 77965 14828 78012
rect 14926 77991 16342 78283
rect 6521 77819 8339 77903
rect 9499 77846 10170 77892
rect 11028 77819 12849 77903
rect 14746 77872 14828 77965
rect 14746 77826 15411 77872
rect 16625 77864 17952 78246
rect 16625 77791 18034 77864
rect 1404 77534 1506 77791
rect 17932 77577 18034 77791
<< metal2 >>
rect 1464 77579 2947 78323
rect 3885 77579 4442 78270
rect 4515 77579 5416 78270
rect 5730 77579 6346 77908
rect 6713 77579 7130 78270
rect 7193 77579 7658 78270
rect 8075 77579 8292 78270
rect 9795 77831 10181 78270
rect 10518 77579 11120 78283
rect 14078 77579 14919 78270
rect 14994 77579 15565 78283
rect 16484 77579 17973 78323
rect 5992 -14 6083 78
rect 8988 -114 9079 -21
rect 9253 -114 9343 -21
rect 9517 -114 9608 -21
rect 9781 -114 9872 -21
rect 10046 -114 10136 -21
rect 10311 -114 10401 -21
rect 11817 -114 11907 -21
rect 12082 -114 12172 -21
rect 12345 -114 12436 -21
rect 12610 -114 12700 -21
rect 12875 -114 12965 -21
rect 13139 -114 13230 -21
rect 13403 -114 13493 -21
rect 13668 -114 13758 -21
<< metal3 >>
rect 48 78138 139 78231
rect 1443 78104 18161 78245
rect 428 77829 517 77922
rect 1443 77807 3714 77948
rect 5730 77815 9434 77908
rect 48 77538 139 77631
rect 9795 77592 9864 77852
rect 15655 77807 18161 77948
rect 18923 77829 19013 77922
rect 0 77236 89 77329
rect 19347 77236 19437 77329
rect 0 76618 89 76711
rect 19347 76618 19437 76711
rect 0 76024 89 76117
rect 19347 76024 19437 76117
rect 0 75406 89 75499
rect 19347 75406 19437 75499
rect 0 74812 89 74905
rect 19347 74812 19437 74905
rect 0 74194 89 74287
rect 19347 74194 19437 74287
rect 0 73600 89 73693
rect 19347 73600 19437 73693
rect 0 72982 89 73075
rect 19347 72982 19437 73075
rect 0 72388 89 72481
rect 19347 72388 19437 72481
rect 0 71770 89 71863
rect 19347 71770 19437 71863
rect 0 71176 89 71269
rect 19347 71176 19437 71269
rect 0 70558 89 70651
rect 19347 70558 19437 70651
rect 0 69964 89 70057
rect 19347 69964 19437 70057
rect 0 69346 89 69439
rect 19347 69346 19437 69439
rect 0 68752 89 68845
rect 19347 68752 19437 68845
rect 0 68134 89 68227
rect 19347 68134 19437 68227
rect 0 67540 89 67633
rect 19347 67540 19437 67633
rect 0 66922 89 67015
rect 19347 66922 19437 67015
rect 0 66328 89 66421
rect 19347 66328 19437 66421
rect 0 65710 89 65803
rect 19347 65710 19437 65803
rect 0 65116 89 65209
rect 19347 65116 19437 65209
rect 0 64498 89 64591
rect 19347 64498 19437 64591
rect 0 63904 89 63997
rect 19347 63904 19437 63997
rect 0 63286 89 63379
rect 19347 63286 19437 63379
rect 0 62692 89 62785
rect 19347 62692 19437 62785
rect 0 62074 89 62167
rect 19347 62074 19437 62167
rect 0 61480 89 61573
rect 19347 61480 19437 61573
rect 0 60862 89 60955
rect 19347 60862 19437 60955
rect 0 60268 89 60361
rect 19347 60268 19437 60361
rect 0 59650 89 59743
rect 19347 59650 19437 59743
rect 0 59056 89 59149
rect 19347 59056 19437 59149
rect 0 58438 89 58531
rect 19347 58438 19437 58531
rect 0 57844 89 57937
rect 19347 57844 19437 57937
rect 0 57226 89 57319
rect 19347 57226 19437 57319
rect 0 56632 89 56725
rect 19347 56632 19437 56725
rect 0 56014 89 56107
rect 19347 56014 19437 56107
rect 0 55420 89 55513
rect 19347 55420 19437 55513
rect 0 54802 89 54895
rect 19347 54802 19437 54895
rect 0 54208 89 54301
rect 19347 54208 19437 54301
rect 0 53590 89 53683
rect 19347 53590 19437 53683
rect 0 52996 89 53089
rect 19347 52996 19437 53089
rect 0 52378 89 52471
rect 19347 52378 19437 52471
rect 0 51784 89 51877
rect 19347 51784 19437 51877
rect 0 51166 89 51259
rect 19347 51166 19437 51259
rect 0 50572 89 50665
rect 19347 50572 19437 50665
rect 0 49954 89 50047
rect 19347 49954 19437 50047
rect 0 49360 89 49453
rect 19347 49360 19437 49453
rect 0 48742 89 48835
rect 19347 48742 19437 48835
rect 0 48148 89 48241
rect 19347 48148 19437 48241
rect 0 47530 89 47623
rect 19347 47530 19437 47623
rect 0 46936 89 47029
rect 19347 46936 19437 47029
rect 0 46318 89 46411
rect 19347 46318 19437 46411
rect 0 45724 89 45817
rect 19347 45724 19437 45817
rect 0 45106 89 45199
rect 19347 45106 19437 45199
rect 0 44512 89 44605
rect 19347 44512 19437 44605
rect 0 43894 89 43987
rect 19347 43894 19437 43987
rect 0 43300 89 43393
rect 19347 43300 19437 43393
rect 0 42682 89 42775
rect 19347 42682 19437 42775
rect 0 42088 89 42181
rect 19347 42088 19437 42181
rect 0 41470 89 41563
rect 19347 41470 19437 41563
rect 0 40876 89 40969
rect 19347 40876 19437 40969
rect 0 40258 89 40351
rect 19347 40258 19437 40351
rect 0 39664 89 39757
rect 19347 39664 19437 39757
rect 0 39046 89 39139
rect 19347 39046 19437 39139
rect 0 38452 89 38545
rect 19347 38452 19437 38545
rect 0 37834 89 37927
rect 19347 37834 19437 37927
rect 0 37240 89 37333
rect 19347 37240 19437 37333
rect 0 36621 89 36714
rect 19347 36622 19437 36715
rect 0 36028 89 36121
rect 19347 36028 19437 36121
rect 0 35410 89 35503
rect 19347 35410 19437 35503
rect 0 34816 89 34909
rect 19347 34816 19437 34909
rect 0 34198 89 34291
rect 19347 34198 19437 34291
rect 0 33604 89 33697
rect 19347 33604 19437 33697
rect 0 32986 89 33079
rect 19347 32986 19437 33079
rect 0 32393 89 32486
rect 19347 32392 19437 32485
rect 0 31774 89 31867
rect 19347 31774 19437 31867
rect 0 31181 89 31274
rect 19347 31180 19437 31273
rect 0 30562 89 30655
rect 19347 30562 19437 30655
rect 0 29969 89 30062
rect 19347 29969 19437 30062
rect 0 29350 89 29443
rect 19347 29351 19437 29444
rect 0 28756 89 28849
rect 19348 28756 19438 28849
rect 0 28138 89 28231
rect 19348 28139 19438 28232
rect 0 27544 89 27637
rect 19348 27545 19438 27638
rect 0 26926 89 27019
rect 19348 26926 19438 27019
rect 0 26333 89 26426
rect 19348 26332 19438 26425
rect 0 25714 89 25807
rect 19348 25714 19438 25807
rect 0 25119 89 25212
rect 19348 25120 19438 25213
rect 0 24502 89 24595
rect 19348 24502 19438 24595
rect 0 23908 89 24001
rect 19348 23908 19438 24001
rect 0 23289 89 23382
rect 19348 23290 19438 23383
rect 0 22696 89 22789
rect 19348 22696 19438 22789
rect 0 22077 89 22170
rect 19348 22077 19438 22170
rect 0 21484 89 21577
rect 19348 21484 19438 21577
rect 0 20865 89 20958
rect 19348 20866 19438 20959
rect 0 20273 89 20366
rect 19348 20272 19438 20365
rect 0 19653 89 19746
rect 19348 19652 19438 19745
rect 0 19059 89 19152
rect 19348 19059 19438 19152
rect 0 18441 89 18534
rect 19348 18443 19438 18536
rect 0 17847 89 17940
rect 19348 17847 19438 17940
rect 0 17231 89 17324
rect 19348 17231 19438 17324
rect 0 16631 89 16724
rect 19348 16635 19438 16728
rect 0 16015 89 16108
rect 19348 16019 19438 16112
rect 0 15423 89 15516
rect 19348 15423 19438 15516
rect 0 14807 89 14900
rect 19348 14807 19438 14900
rect 0 14211 89 14304
rect 19348 14211 19438 14304
rect 0 13595 89 13688
rect 19348 13595 19438 13688
rect 0 12999 89 13092
rect 19348 12999 19438 13092
rect 0 12383 89 12476
rect 19348 12383 19438 12476
rect 0 11787 89 11880
rect 19348 11787 19438 11880
rect 0 11171 89 11264
rect 19348 11171 19438 11264
rect 0 10575 89 10668
rect 19348 10575 19438 10668
rect 0 9959 89 10052
rect 19348 9959 19438 10052
rect 0 9363 89 9456
rect 19348 9363 19438 9456
rect 0 8747 89 8840
rect 19348 8747 19438 8840
rect 0 8150 89 8243
rect 19348 8151 19438 8244
rect 0 7534 89 7627
rect 19348 7535 19438 7628
rect 0 6939 89 7032
rect 19348 6939 19438 7032
rect 0 6323 89 6416
rect 19348 6323 19438 6416
rect 0 5727 89 5820
rect 19348 5727 19438 5820
rect 0 5111 89 5204
rect 19348 5111 19438 5204
rect 0 4515 89 4608
rect 19348 4515 19438 4608
rect 0 3899 89 3992
rect 19348 3899 19438 3992
rect 0 3301 89 3394
rect 19348 3301 19438 3394
rect 0 2685 89 2778
rect 19348 2685 19438 2778
rect 0 2091 89 2184
rect 19348 2091 19438 2184
rect 0 1475 89 1568
rect 19348 1475 19438 1568
rect 0 880 89 973
rect 19348 881 19438 974
rect 0 263 89 356
rect 19348 265 19438 358
use M1_NACTIVE_02_3v1024x8m81  M1_NACTIVE_02_3v1024x8m81_0
timestamp 1764525316
transform 1 0 9844 0 1 78241
box -54 -56 607 56
use M1_NWELL_01_3v1024x8m81  M1_NWELL_01_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1540 0 1 78190
box -154 -501 1372 159
use M1_NWELL_01_3v1024x8m81  M1_NWELL_01_3v1024x8m81_1
timestamp 1764525316
transform -1 0 17897 0 1 78190
box -154 -501 1372 159
use M1_PACTIVE$10_3v1024x8m81  M1_PACTIVE$10_3v1024x8m81_0
timestamp 1764525316
transform 1 0 8024 0 1 78241
box -54 -56 1271 56
use M1_PACTIVE$10_3v1024x8m81  M1_PACTIVE$10_3v1024x8m81_1
timestamp 1764525316
transform 1 0 3073 0 1 78241
box -54 -56 1271 56
use M1_PACTIVE$10_3v1024x8m81  M1_PACTIVE$10_3v1024x8m81_2
timestamp 1764525316
transform 1 0 15032 0 1 78241
box -54 -56 1271 56
use M1_PACTIVE$11_3v1024x8m81  M1_PACTIVE$11_3v1024x8m81_0
timestamp 1764525316
transform 1 0 11102 0 1 78241
box -54 -56 275 56
use M1_POLY2$$204150828_3v1024x8m81  M1_POLY2$$204150828_3v1024x8m81_0
timestamp 1764525316
transform 1 0 6561 0 1 77988
box -46 -122 46 122
use M1_POLY24310591302019_3v1024x8m81  M1_POLY24310591302019_3v1024x8m81_0
timestamp 1764525316
transform 1 0 8428 0 1 77962
box -36 -80 36 78
use M1_POLY24310591302019_3v1024x8m81  M1_POLY24310591302019_3v1024x8m81_1
timestamp 1764525316
transform 0 -1 9598 1 0 78195
box -36 -80 36 78
use M1_POLY24310591302019_3v1024x8m81  M1_POLY24310591302019_3v1024x8m81_2
timestamp 1764525316
transform 1 0 10937 0 1 77990
box -36 -80 36 78
use M1_POLY24310591302019_3v1024x8m81  M1_POLY24310591302019_3v1024x8m81_3
timestamp 1764525316
transform 1 0 12819 0 1 77990
box -36 -80 36 78
use M1_POLY24310591302031_3v1024x8m81  M1_POLY24310591302031_3v1024x8m81_0
timestamp 1764525316
transform 1 0 10789 0 1 78228
box -36 -36 36 36
use M2_M1$$201262124_3v1024x8m81  M2_M1$$201262124_3v1024x8m81_0
timestamp 1764525316
transform 1 0 9590 0 1 78193
box -119 -46 119 46
use M2_M1$$204138540_3v1024x8m81  M2_M1$$204138540_3v1024x8m81_0
timestamp 1764525316
transform 1 0 7281 0 1 78023
box -45 -46 340 46
use M2_M1$$204138540_3v1024x8m81  M2_M1$$204138540_3v1024x8m81_1
timestamp 1764525316
transform 1 0 9841 0 1 78236
box -45 -46 340 46
use M2_M1$$204139564_3v1024x8m81  M2_M1$$204139564_3v1024x8m81_0
timestamp 1764525316
transform 1 0 8120 0 1 78203
box -45 -198 171 46
use M2_M1$$204140588_3v1024x8m81  M2_M1$$204140588_3v1024x8m81_0
timestamp 1764525316
transform 1 0 8651 0 1 77861
box -45 -46 783 46
use M2_M1$$204141612_3v1024x8m81  M2_M1$$204141612_3v1024x8m81_0
timestamp 1764525316
transform 1 0 10588 0 1 78236
box -45 -46 487 46
use M2_M1$$204141612_3v1024x8m81  M2_M1$$204141612_3v1024x8m81_1
timestamp 1764525316
transform 1 0 14123 0 1 78186
box -45 -46 487 46
use M2_M1$$204141612_3v1024x8m81  M2_M1$$204141612_3v1024x8m81_2
timestamp 1764525316
transform 1 0 14123 0 1 77861
box -45 -46 487 46
use M2_M1$$204220460_3v1024x8m81  M2_M1$$204220460_3v1024x8m81_0
timestamp 1764525316
transform 1 0 3079 0 1 77863
box -45 -46 635 46
use M2_M1$$204220460_3v1024x8m81  M2_M1$$204220460_3v1024x8m81_1
timestamp 1764525316
transform 1 0 4754 0 1 78151
box -45 -46 635 46
use M2_M1$$204220460_3v1024x8m81  M2_M1$$204220460_3v1024x8m81_2
timestamp 1764525316
transform 1 0 4754 0 1 77826
box -45 -46 635 46
use M2_M1$$204220460_3v1024x8m81  M2_M1$$204220460_3v1024x8m81_3
timestamp 1764525316
transform 1 0 15701 0 1 77861
box -45 -46 635 46
use M2_M1$$204221484_3v1024x8m81  M2_M1$$204221484_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1509 0 1 78200
box -45 -351 1225 46
use M2_M1$$204221484_3v1024x8m81  M2_M1$$204221484_3v1024x8m81_1
timestamp 1764525316
transform -1 0 17928 0 1 78200
box -45 -351 1225 46
use M2_M1$$204222508_3v1024x8m81  M2_M1$$204222508_3v1024x8m81_0
timestamp 1764525316
transform 1 0 3947 0 1 78200
box -45 -198 487 46
use M2_M1$$204222508_3v1024x8m81  M2_M1$$204222508_3v1024x8m81_1
timestamp 1764525316
transform 1 0 15040 0 1 78200
box -45 -198 487 46
use M3_M2$$204142636_3v1024x8m81  M3_M2$$204142636_3v1024x8m81_0
timestamp 1764525316
transform 1 0 3947 0 1 78200
box -44 -46 487 46
use M3_M2$$204142636_3v1024x8m81  M3_M2$$204142636_3v1024x8m81_1
timestamp 1764525316
transform 1 0 5775 0 1 77861
box -44 -46 487 46
use M3_M2$$204142636_3v1024x8m81  M3_M2$$204142636_3v1024x8m81_3
timestamp 1764525316
transform 1 0 15040 0 1 78200
box -44 -46 487 46
use M3_M2$$204143660_3v1024x8m81  M3_M2$$204143660_3v1024x8m81_0
timestamp 1764525316
transform 1 0 8120 0 1 78200
box -45 -46 171 46
use M3_M2$$204144684_3v1024x8m81  M3_M2$$204144684_3v1024x8m81_0
timestamp 1764525316
transform 1 0 3079 0 1 77863
box -45 -46 635 46
use M3_M2$$204144684_3v1024x8m81  M3_M2$$204144684_3v1024x8m81_1
timestamp 1764525316
transform 1 0 15701 0 1 77861
box -45 -46 635 46
use M3_M2$$204145708_3v1024x8m81  M3_M2$$204145708_3v1024x8m81_0
timestamp 1764525316
transform 1 0 8651 0 1 77861
box -45 -46 783 46
use M3_M2$$204146732_3v1024x8m81  M3_M2$$204146732_3v1024x8m81_0
timestamp 1764525316
transform 1 0 9841 0 1 77857
box -45 -46 340 46
use nmos_1p2_01_R270_3v1024x8m81  nmos_1p2_01_R270_3v1024x8m81_0
timestamp 1764525316
transform 0 -1 9522 -1 0 77963
box -102 -44 130 659
use nmos_1p2_02_R90_3v1024x8m81  nmos_1p2_02_R90_3v1024x8m81_0
timestamp 1764525316
transform 0 -1 4442 1 0 77922
box -102 -44 130 987
use nmos_5p04310591302099_3v1024x8m81  nmos_5p04310591302099_3v1024x8m81_0
timestamp 1764525316
transform 0 -1 16342 1 0 77900
box -88 -44 144 987
use nmos_5p043105913020111_3v1024x8m81  nmos_5p043105913020111_3v1024x8m81_0
timestamp 1764525316
transform 0 -1 8339 1 0 77900
box -88 -44 144 291
use nmos_5p043105913020111_3v1024x8m81  nmos_5p043105913020111_3v1024x8m81_1
timestamp 1764525316
transform 0 -1 11398 1 0 77900
box -88 -44 144 291
use pmos_1p2_01_R90_3v1024x8m81  pmos_1p2_01_R90_3v1024x8m81_0
timestamp 1764525316
transform 0 -1 7702 1 0 77922
box -188 -86 216 701
use pmos_1p2_02_R90_3v1024x8m81  pmos_1p2_02_R90_3v1024x8m81_0
timestamp 1764525316
transform 0 -1 6471 1 0 77922
box -216 -86 348 1264
use pmos_1p2_02_R90_3v1024x8m81  pmos_1p2_02_R90_3v1024x8m81_1
timestamp 1764525316
transform 0 -1 14665 1 0 77922
box -216 -86 348 1264
use pmos_5p043105913020101_3v1024x8m81  pmos_5p043105913020101_3v1024x8m81_0
timestamp 1764525316
transform 0 -1 12581 1 0 77900
box -174 -86 230 701
use pmos_5p043105913020101_3v1024x8m81  pmos_5p043105913020101_3v1024x8m81_1
timestamp 1764525316
transform 0 -1 10712 1 0 77900
box -174 -86 230 701
use pmoscap_L1_W2_R270_3v1024x8m81  pmoscap_L1_W2_R270_3v1024x8m81_0
timestamp 1764692000
transform 0 -1 1542 -1 0 78230
box -88 -189 771 1517
use pmoscap_L1_W2_R270_3v1024x8m81  pmoscap_L1_W2_R270_3v1024x8m81_1
timestamp 1764692000
transform 0 1 17896 -1 0 78230
box -88 -189 771 1517
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_0
timestamp 1764525316
transform 0 1 17896 -1 0 10822
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_1
timestamp 1764525316
transform 0 1 17896 -1 0 9610
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_2
timestamp 1764525316
transform 0 1 17896 -1 0 8398
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_3
timestamp 1764525316
transform 0 1 17896 -1 0 7186
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_4
timestamp 1764525316
transform 0 1 17896 -1 0 5974
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_5
timestamp 1764525316
transform 0 1 17896 -1 0 4762
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_6
timestamp 1764525316
transform 0 1 17896 -1 0 3550
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_7
timestamp 1764525316
transform 0 1 17896 -1 0 2338
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_8
timestamp 1764525316
transform 0 1 17896 -1 0 1126
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_9
timestamp 1764525316
transform 0 1 17896 -1 0 19306
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_10
timestamp 1764525316
transform 0 1 17896 -1 0 18094
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_11
timestamp 1764525316
transform 0 1 17896 -1 0 16882
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_12
timestamp 1764525316
transform 0 1 17896 -1 0 15670
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_13
timestamp 1764525316
transform 0 1 17896 -1 0 14458
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_14
timestamp 1764525316
transform 0 1 17896 -1 0 13246
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_15
timestamp 1764525316
transform 0 1 17896 -1 0 12034
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_16
timestamp 1764525316
transform 0 -1 1542 -1 0 10822
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_17
timestamp 1764525316
transform 0 -1 1542 -1 0 9610
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_18
timestamp 1764525316
transform 0 -1 1542 -1 0 8398
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_19
timestamp 1764525316
transform 0 -1 1542 -1 0 7186
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_20
timestamp 1764525316
transform 0 -1 1542 -1 0 5974
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_21
timestamp 1764525316
transform 0 -1 1542 -1 0 4762
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_22
timestamp 1764525316
transform 0 -1 1542 -1 0 3550
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_23
timestamp 1764525316
transform 0 -1 1542 -1 0 2338
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_24
timestamp 1764525316
transform 0 -1 1542 -1 0 1126
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_25
timestamp 1764525316
transform 0 -1 1542 -1 0 19306
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_26
timestamp 1764525316
transform 0 -1 1542 -1 0 18094
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_27
timestamp 1764525316
transform 0 -1 1542 -1 0 16882
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_28
timestamp 1764525316
transform 0 -1 1542 -1 0 15670
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_29
timestamp 1764525316
transform 0 -1 1542 -1 0 14458
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_30
timestamp 1764525316
transform 0 -1 1542 -1 0 13246
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_31
timestamp 1764525316
transform 0 -1 1542 -1 0 12034
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_32
timestamp 1764525316
transform 0 -1 1542 -1 0 38698
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_33
timestamp 1764525316
transform 0 -1 1542 -1 0 37486
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_34
timestamp 1764525316
transform 0 -1 1542 -1 0 36274
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_35
timestamp 1764525316
transform 0 -1 1542 -1 0 35062
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_36
timestamp 1764525316
transform 0 -1 1542 -1 0 33850
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_37
timestamp 1764525316
transform 0 -1 1542 -1 0 32638
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_38
timestamp 1764525316
transform 0 -1 1542 -1 0 31426
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_39
timestamp 1764525316
transform 0 -1 1542 -1 0 30214
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_40
timestamp 1764525316
transform 0 -1 1542 -1 0 29002
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_41
timestamp 1764525316
transform 0 -1 1542 -1 0 27790
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_42
timestamp 1764525316
transform 0 -1 1542 -1 0 26578
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_43
timestamp 1764525316
transform 0 -1 1542 -1 0 25366
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_44
timestamp 1764525316
transform 0 -1 1542 -1 0 24154
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_45
timestamp 1764525316
transform 0 -1 1542 -1 0 22942
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_46
timestamp 1764525316
transform 0 -1 1542 -1 0 21730
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_47
timestamp 1764525316
transform 0 1 17896 -1 0 38698
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_48
timestamp 1764525316
transform 0 1 17896 -1 0 37486
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_49
timestamp 1764525316
transform 0 1 17896 -1 0 36274
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_50
timestamp 1764525316
transform 0 1 17896 -1 0 35062
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_51
timestamp 1764525316
transform 0 1 17896 -1 0 33850
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_52
timestamp 1764525316
transform 0 1 17896 -1 0 32638
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_53
timestamp 1764525316
transform 0 1 17896 -1 0 31426
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_54
timestamp 1764525316
transform 0 1 17896 -1 0 30214
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_55
timestamp 1764525316
transform 0 1 17896 -1 0 29002
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_56
timestamp 1764525316
transform 0 1 17896 -1 0 27790
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_57
timestamp 1764525316
transform 0 1 17896 -1 0 26578
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_58
timestamp 1764525316
transform 0 1 17896 -1 0 25366
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_59
timestamp 1764525316
transform 0 1 17896 -1 0 24154
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_60
timestamp 1764525316
transform 0 1 17896 -1 0 22942
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_61
timestamp 1764525316
transform 0 1 17896 -1 0 21730
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_62
timestamp 1764525316
transform 0 -1 1542 -1 0 20518
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_63
timestamp 1764525316
transform 0 1 17896 -1 0 20518
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_64
timestamp 1764525316
transform 0 -1 1542 -1 0 39910
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_65
timestamp 1764525316
transform 0 1 17896 -1 0 39910
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_66
timestamp 1764525316
transform 0 -1 1542 -1 0 41122
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_67
timestamp 1764525316
transform 0 1 17896 -1 0 41122
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_68
timestamp 1764525316
transform 0 -1 1542 -1 0 42334
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_69
timestamp 1764525316
transform 0 1 17896 -1 0 42334
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_70
timestamp 1764525316
transform 0 -1 1542 -1 0 43546
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_71
timestamp 1764525316
transform 0 1 17896 -1 0 43546
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_72
timestamp 1764525316
transform 0 -1 1542 -1 0 44758
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_73
timestamp 1764525316
transform 0 1 17896 -1 0 44758
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_74
timestamp 1764525316
transform 0 -1 1542 -1 0 45970
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_75
timestamp 1764525316
transform 0 1 17896 -1 0 45970
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_76
timestamp 1764525316
transform 0 -1 1542 -1 0 47182
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_77
timestamp 1764525316
transform 0 1 17896 -1 0 47182
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_78
timestamp 1764525316
transform 0 -1 1542 -1 0 48394
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_79
timestamp 1764525316
transform 0 1 17896 -1 0 48394
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_80
timestamp 1764525316
transform 0 -1 1542 -1 0 49606
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_81
timestamp 1764525316
transform 0 1 17896 -1 0 49606
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_82
timestamp 1764525316
transform 0 -1 1542 -1 0 50818
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_83
timestamp 1764525316
transform 0 1 17896 -1 0 50818
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_84
timestamp 1764525316
transform 0 -1 1542 -1 0 52030
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_85
timestamp 1764525316
transform 0 1 17896 -1 0 52030
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_86
timestamp 1764525316
transform 0 -1 1542 -1 0 53242
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_87
timestamp 1764525316
transform 0 1 17896 -1 0 53242
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_88
timestamp 1764525316
transform 0 -1 1542 -1 0 54454
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_89
timestamp 1764525316
transform 0 1 17896 -1 0 54454
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_90
timestamp 1764525316
transform 0 -1 1542 -1 0 55666
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_91
timestamp 1764525316
transform 0 1 17896 -1 0 55666
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_92
timestamp 1764525316
transform 0 -1 1542 -1 0 56878
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_93
timestamp 1764525316
transform 0 1 17896 -1 0 56878
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_94
timestamp 1764525316
transform 0 -1 1542 -1 0 58090
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_95
timestamp 1764525316
transform 0 1 17896 -1 0 58090
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_96
timestamp 1764525316
transform 0 -1 1542 -1 0 59302
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_97
timestamp 1764525316
transform 0 1 17896 -1 0 59302
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_98
timestamp 1764525316
transform 0 -1 1542 -1 0 60514
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_99
timestamp 1764525316
transform 0 1 17896 -1 0 60514
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_100
timestamp 1764525316
transform 0 -1 1542 -1 0 61726
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_101
timestamp 1764525316
transform 0 1 17896 -1 0 61726
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_102
timestamp 1764525316
transform 0 -1 1542 -1 0 62938
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_103
timestamp 1764525316
transform 0 1 17896 -1 0 62938
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_104
timestamp 1764525316
transform 0 -1 1542 -1 0 64150
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_105
timestamp 1764525316
transform 0 1 17896 -1 0 64150
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_106
timestamp 1764525316
transform 0 -1 1542 -1 0 65362
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_107
timestamp 1764525316
transform 0 1 17896 -1 0 65362
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_108
timestamp 1764525316
transform 0 -1 1542 -1 0 66574
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_109
timestamp 1764525316
transform 0 1 17896 -1 0 66574
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_110
timestamp 1764525316
transform 0 -1 1542 -1 0 67786
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_111
timestamp 1764525316
transform 0 1 17896 -1 0 67786
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_112
timestamp 1764525316
transform 0 -1 1542 -1 0 68998
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_113
timestamp 1764525316
transform 0 1 17896 -1 0 68998
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_114
timestamp 1764525316
transform 0 -1 1542 -1 0 70210
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_115
timestamp 1764525316
transform 0 1 17896 -1 0 70210
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_116
timestamp 1764525316
transform 0 -1 1542 -1 0 71422
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_117
timestamp 1764525316
transform 0 1 17896 -1 0 71422
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_118
timestamp 1764525316
transform 0 -1 1542 -1 0 72634
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_119
timestamp 1764525316
transform 0 1 17896 -1 0 72634
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_120
timestamp 1764525316
transform 0 -1 1542 -1 0 73846
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_121
timestamp 1764525316
transform 0 1 17896 -1 0 73846
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_122
timestamp 1764525316
transform 0 -1 1542 -1 0 75058
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_123
timestamp 1764525316
transform 0 1 17896 -1 0 75058
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_124
timestamp 1764525316
transform 0 -1 1542 -1 0 76270
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_125
timestamp 1764525316
transform 0 1 17896 -1 0 76270
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_126
timestamp 1764525316
transform 0 -1 1542 -1 0 77482
box -226 -219 1235 3808
use pmoscap_R270_3v1024x8m81  pmoscap_R270_3v1024x8m81_127
timestamp 1764525316
transform 0 1 17896 -1 0 77482
box -226 -219 1235 3808
use xdec32_3v1024x8m81  xdec32_3v1024x8m81_0
timestamp 1764692000
transform 1 0 1208 0 1 0
box 230 -159 16952 19575
use xdec32_468_3v1024x8m81  xdec32_468_3v1024x8m81_0
timestamp 1764692000
transform 1 0 1208 0 1 19392
box 230 -159 16952 19575
use xdec64_3v1024x8m81  xdec64_3v1024x8m81_0
timestamp 1765483240
transform 1 0 1208 0 1 38784
box 230 -159 16952 19575
use xdec64_468_3v1024x8m81  xdec64_468_3v1024x8m81_0
timestamp 1765483240
transform 1 0 1208 0 1 58176
box 230 -159 16952 19575
<< labels >>
rlabel metal2 s 10355 -67 10355 -67 4 xb[0]
port 133 nsew
rlabel metal2 s 10091 -67 10091 -67 4 xb[1]
port 134 nsew
rlabel metal2 s 9827 -67 9827 -67 4 xb[2]
port 135 nsew
rlabel metal2 s 9562 -67 9562 -67 4 xb[3]
port 136 nsew
rlabel metal2 s 11862 -67 11862 -67 4 xa[7]
port 137 nsew
rlabel metal2 s 12126 -67 12126 -67 4 xa[6]
port 138 nsew
rlabel metal2 s 12391 -67 12391 -67 4 xa[5]
port 139 nsew
rlabel metal2 s 12656 -67 12656 -67 4 xa[4]
port 140 nsew
rlabel metal2 s 13713 -67 13713 -67 4 xa[0]
port 141 nsew
rlabel metal2 s 6038 31 6038 31 4 men
port 142 nsew
rlabel metal2 s 12919 -67 12919 -67 4 xa[3]
port 143 nsew
rlabel metal2 s 13184 -67 13184 -67 4 xa[2]
port 144 nsew
rlabel metal2 s 13449 -67 13449 -67 4 xa[1]
port 145 nsew
rlabel metal2 s 9298 -67 9298 -67 4 xc[0]
port 146 nsew
rlabel metal2 s 9034 -67 9034 -67 4 xc[1]
port 147 nsew
rlabel metal3 s 44 927 44 927 4 LWL[1]
port 91 nsew
rlabel metal3 s 44 310 44 310 4 LWL[0]
port 92 nsew
rlabel metal3 s 44 1522 44 1522 4 LWL[2]
port 90 nsew
rlabel metal3 s 44 2138 44 2138 4 LWL[3]
port 89 nsew
rlabel metal3 s 44 2732 44 2732 4 LWL[4]
port 88 nsew
rlabel metal3 s 44 3348 44 3348 4 LWL[5]
port 87 nsew
rlabel metal3 s 44 3946 44 3946 4 LWL[6]
port 95 nsew
rlabel metal3 s 44 4562 44 4562 4 LWL[7]
port 97 nsew
rlabel metal3 s 44 5158 44 5158 4 LWL[8]
port 93 nsew
rlabel metal3 s 44 5774 44 5774 4 LWL[9]
port 94 nsew
rlabel metal3 s 44 6370 44 6370 4 LWL[10]
port 78 nsew
rlabel metal3 s 44 6986 44 6986 4 LWL[11]
port 79 nsew
rlabel metal3 s 44 7581 44 7581 4 LWL[12]
port 80 nsew
rlabel metal3 s 44 8197 44 8197 4 LWL[13]
port 81 nsew
rlabel metal3 s 44 8794 44 8794 4 LWL[14]
port 82 nsew
rlabel metal3 s 44 9410 44 9410 4 LWL[15]
port 83 nsew
rlabel metal3 s 44 10006 44 10006 4 LWL[16]
port 84 nsew
rlabel metal3 s 44 10622 44 10622 4 LWL[17]
port 85 nsew
rlabel metal3 s 44 11218 44 11218 4 LWL[18]
port 86 nsew
rlabel metal3 s 44 11834 44 11834 4 LWL[19]
port 68 nsew
rlabel metal3 s 44 13046 44 13046 4 LWL[21]
port 70 nsew
rlabel metal3 s 44 12430 44 12430 4 LWL[20]
port 69 nsew
rlabel metal3 s 44 13642 44 13642 4 LWL[22]
port 71 nsew
rlabel metal3 s 44 14258 44 14258 4 LWL[23]
port 72 nsew
rlabel metal3 s 44 14854 44 14854 4 LWL[24]
port 73 nsew
rlabel metal3 s 44 15470 44 15470 4 LWL[25]
port 74 nsew
rlabel metal3 s 44 16062 44 16062 4 LWL[26]
port 75 nsew
rlabel metal3 s 44 16678 44 16678 4 LWL[27]
port 76 nsew
rlabel metal3 s 44 18488 44 18488 4 LWL[30]
port 99 nsew
rlabel metal3 s 44 17894 44 17894 4 LWL[29]
port 98 nsew
rlabel metal3 s 44 17278 44 17278 4 LWL[28]
port 77 nsew
rlabel metal3 s 44 19106 44 19106 4 LWL[31]
port 67 nsew
rlabel metal3 s 44 21531 44 21531 4 LWL[35]
port 61 nsew
rlabel metal3 s 44 20912 44 20912 4 LWL[34]
port 62 nsew
rlabel metal3 s 44 20320 44 20320 4 LWL[33]
port 63 nsew
rlabel metal3 s 44 19700 44 19700 4 LWL[32]
port 96 nsew
rlabel metal3 s 44 22124 44 22124 4 LWL[36]
port 60 nsew
rlabel metal3 s 44 22743 44 22743 4 LWL[37]
port 59 nsew
rlabel metal3 s 44 23336 44 23336 4 LWL[38]
port 58 nsew
rlabel metal3 s 44 23955 44 23955 4 LWL[39]
port 57 nsew
rlabel metal3 s 44 24549 44 24549 4 LWL[40]
port 56 nsew
rlabel metal3 s 44 25166 44 25166 4 LWL[41]
port 55 nsew
rlabel metal3 s 44 25761 44 25761 4 LWL[42]
port 54 nsew
rlabel metal3 s 44 26380 44 26380 4 LWL[43]
port 53 nsew
rlabel metal3 s 44 26973 44 26973 4 LWL[44]
port 52 nsew
rlabel metal3 s 44 27591 44 27591 4 LWL[45]
port 51 nsew
rlabel metal3 s 44 28185 44 28185 4 LWL[46]
port 50 nsew
rlabel metal3 s 44 28803 44 28803 4 LWL[47]
port 49 nsew
rlabel metal3 s 44 29397 44 29397 4 LWL[48]
port 48 nsew
rlabel metal3 s 44 30016 44 30016 4 LWL[49]
port 47 nsew
rlabel metal3 s 44 30609 44 30609 4 LWL[50]
port 46 nsew
rlabel metal3 s 44 31228 44 31228 4 LWL[51]
port 45 nsew
rlabel metal3 s 44 31821 44 31821 4 LWL[52]
port 44 nsew
rlabel metal3 s 44 32440 44 32440 4 LWL[53]
port 43 nsew
rlabel metal3 s 44 33033 44 33033 4 LWL[54]
port 42 nsew
rlabel metal3 s 44 33651 44 33651 4 LWL[55]
port 41 nsew
rlabel metal3 s 44 34245 44 34245 4 LWL[56]
port 40 nsew
rlabel metal3 s 44 34863 44 34863 4 LWL[57]
port 39 nsew
rlabel metal3 s 44 35457 44 35457 4 LWL[58]
port 38 nsew
rlabel metal3 s 44 36075 44 36075 4 LWL[59]
port 37 nsew
rlabel metal3 s 44 36668 44 36668 4 LWL[60]
port 36 nsew
rlabel metal3 s 35 38506 35 38506 4 LWL[63]
port 33 nsew
rlabel metal3 s 19393 928 19393 928 4 RWL[1]
port 116 nsew
rlabel metal3 s 19393 312 19393 312 4 RWL[0]
port 115 nsew
rlabel metal3 s 19393 1522 19393 1522 4 RWL[2]
port 114 nsew
rlabel metal3 s 19393 2138 19393 2138 4 RWL[3]
port 117 nsew
rlabel metal3 s 19393 2732 19393 2732 4 RWL[4]
port 113 nsew
rlabel metal3 s 19393 3348 19393 3348 4 RWL[5]
port 118 nsew
rlabel metal3 s 19393 3946 19393 3946 4 RWL[6]
port 112 nsew
rlabel metal3 s 19393 4562 19393 4562 4 RWL[7]
port 119 nsew
rlabel metal3 s 19393 5158 19393 5158 4 RWL[8]
port 120 nsew
rlabel metal3 s 19393 5774 19393 5774 4 RWL[9]
port 121 nsew
rlabel metal3 s 19393 6370 19393 6370 4 RWL[10]
port 122 nsew
rlabel metal3 s 19393 6986 19393 6986 4 RWL[11]
port 123 nsew
rlabel metal3 s 19393 7582 19393 7582 4 RWL[12]
port 124 nsew
rlabel metal3 s 19393 8198 19393 8198 4 RWL[13]
port 125 nsew
rlabel metal3 s 19393 8794 19393 8794 4 RWL[14]
port 126 nsew
rlabel metal3 s 19393 9410 19393 9410 4 RWL[15]
port 127 nsew
rlabel metal3 s 19393 10006 19393 10006 4 RWL[16]
port 128 nsew
rlabel metal3 s 19393 10622 19393 10622 4 RWL[17]
port 129 nsew
rlabel metal3 s 19393 11218 19393 11218 4 RWL[18]
port 130 nsew
rlabel metal3 s 19393 11834 19393 11834 4 RWL[19]
port 131 nsew
rlabel metal3 s 19393 13046 19393 13046 4 RWL[21]
port 111 nsew
rlabel metal3 s 19393 12430 19393 12430 4 RWL[20]
port 132 nsew
rlabel metal3 s 19393 13642 19393 13642 4 RWL[22]
port 110 nsew
rlabel metal3 s 19393 14258 19393 14258 4 RWL[23]
port 109 nsew
rlabel metal3 s 19393 15470 19393 15470 4 RWL[25]
port 107 nsew
rlabel metal3 s 19393 14854 19393 14854 4 RWL[24]
port 108 nsew
rlabel metal3 s 19393 16682 19393 16682 4 RWL[27]
port 105 nsew
rlabel metal3 s 19393 16066 19393 16066 4 RWL[26]
port 106 nsew
rlabel metal3 s 19393 17894 19393 17894 4 RWL[29]
port 103 nsew
rlabel metal3 s 19393 17278 19393 17278 4 RWL[28]
port 104 nsew
rlabel metal3 s 19393 19106 19393 19106 4 RWL[31]
port 101 nsew
rlabel metal3 s 19393 18490 19393 18490 4 RWL[30]
port 102 nsew
rlabel metal3 s 19393 19699 19393 19699 4 RWL[32]
port 100 nsew
rlabel metal3 s 19393 20319 19393 20319 4 RWL[33]
port 2 nsew
rlabel metal3 s 19393 20913 19393 20913 4 RWL[34]
port 3 nsew
rlabel metal3 s 19393 21531 19393 21531 4 RWL[35]
port 4 nsew
rlabel metal3 s 19393 22124 19393 22124 4 RWL[36]
port 5 nsew
rlabel metal3 s 19393 22743 19393 22743 4 RWL[37]
port 6 nsew
rlabel metal3 s 19393 23337 19393 23337 4 RWL[38]
port 7 nsew
rlabel metal3 s 19393 23955 19393 23955 4 RWL[39]
port 8 nsew
rlabel metal3 s 19393 24549 19393 24549 4 RWL[40]
port 9 nsew
rlabel metal3 s 19393 25167 19393 25167 4 RWL[41]
port 10 nsew
rlabel metal3 s 19393 25761 19393 25761 4 RWL[42]
port 11 nsew
rlabel metal3 s 19393 26379 19393 26379 4 RWL[43]
port 12 nsew
rlabel metal3 s 19393 26973 19393 26973 4 RWL[44]
port 13 nsew
rlabel metal3 s 19393 27592 19393 27592 4 RWL[45]
port 14 nsew
rlabel metal3 s 19393 28186 19393 28186 4 RWL[46]
port 15 nsew
rlabel metal3 s 19393 28803 19393 28803 4 RWL[47]
port 16 nsew
rlabel metal3 s 19392 29398 19392 29398 4 RWL[48]
port 17 nsew
rlabel metal3 s 19392 30016 19392 30016 4 RWL[49]
port 18 nsew
rlabel metal3 s 19392 30609 19392 30609 4 RWL[50]
port 19 nsew
rlabel metal3 s 19392 31227 19392 31227 4 RWL[51]
port 20 nsew
rlabel metal3 s 19392 31821 19392 31821 4 RWL[52]
port 21 nsew
rlabel metal3 s 19392 32439 19392 32439 4 RWL[53]
port 22 nsew
rlabel metal3 s 19392 33033 19392 33033 4 RWL[54]
port 23 nsew
rlabel metal3 s 19392 33651 19392 33651 4 RWL[55]
port 24 nsew
rlabel metal3 s 19392 34245 19392 34245 4 RWL[56]
port 25 nsew
rlabel metal3 s 19392 34863 19392 34863 4 RWL[57]
port 26 nsew
rlabel metal3 s 19392 35457 19392 35457 4 RWL[58]
port 27 nsew
rlabel metal3 s 19392 36075 19392 36075 4 RWL[59]
port 28 nsew
rlabel metal3 s 19392 36669 19392 36669 4 RWL[60]
port 29 nsew
rlabel metal3 s 19392 37287 19392 37287 4 RWL[61]
port 30 nsew
rlabel metal3 s 19392 37881 19392 37881 4 RWL[62]
port 31 nsew
rlabel metal3 s 19392 38499 19392 38499 4 RWL[63]
port 32 nsew
rlabel metal3 s 93 77585 93 77585 4 vdd
port 65 nsew
rlabel metal3 s 472 77876 472 77876 4 DLWL
port 66 nsew
rlabel metal3 s 18968 77876 18968 77876 4 DRWL
port 1 nsew
rlabel metal3 s 93 78185 93 78185 4 vss
port 64 nsew
rlabel metal3 s 44 37297 44 37297 4 LWL[61]
port 35 nsew
rlabel metal3 s 44 37891 44 37891 4 LWL[62]
port 34 nsew
rlabel metal3 19390 39092 19390 39092 0 RWL[64]
port 148 nsew
rlabel metal3 19390 39714 19390 39714 0 RWL[65]
port 149 nsew
rlabel metal3 19390 40304 19390 40304 0 RWL[66]
port 150 nsew
rlabel metal3 19390 40926 19390 40926 0 RWL[67]
port 151 nsew
rlabel metal3 19390 41516 19390 41516 0 RWL[68]
port 152 nsew
rlabel metal3 19390 42138 19390 42138 0 RWL[69]
port 153 nsew
rlabel metal3 19390 42728 19390 42728 0 RWL[70]
port 154 nsew
rlabel metal3 19390 43350 19390 43350 0 RWL[71]
port 155 nsew
rlabel metal3 19390 43940 19390 43940 0 RWL[72]
port 156 nsew
rlabel metal3 19390 44562 19390 44562 0 RWL[73]
port 157 nsew
rlabel metal3 19390 45152 19390 45152 0 RWL[74]
port 158 nsew
rlabel metal3 19390 45774 19390 45774 0 RWL[75]
port 159 nsew
rlabel metal3 19390 46364 19390 46364 0 RWL[76]
port 160 nsew
rlabel metal3 19390 46986 19390 46986 0 RWL[77]
port 161 nsew
rlabel metal3 19390 47576 19390 47576 0 RWL[78]
port 162 nsew
rlabel metal3 19390 48198 19390 48198 0 RWL[79]
port 163 nsew
rlabel metal3 19390 48788 19390 48788 0 RWL[80]
port 164 nsew
rlabel metal3 19390 49410 19390 49410 0 RWL[81]
port 165 nsew
rlabel metal3 19390 50000 19390 50000 0 RWL[82]
port 166 nsew
rlabel metal3 19390 50622 19390 50622 0 RWL[83]
port 167 nsew
rlabel metal3 19390 51212 19390 51212 0 RWL[84]
port 168 nsew
rlabel metal3 19390 51834 19390 51834 0 RWL[85]
port 169 nsew
rlabel metal3 19390 52424 19390 52424 0 RWL[86]
port 170 nsew
rlabel metal3 19390 53046 19390 53046 0 RWL[87]
port 171 nsew
rlabel metal3 19390 53636 19390 53636 0 RWL[88]
port 172 nsew
rlabel metal3 19390 54258 19390 54258 0 RWL[89]
port 173 nsew
rlabel metal3 19390 54848 19390 54848 0 RWL[90]
port 174 nsew
rlabel metal3 19390 55470 19390 55470 0 RWL[91]
port 175 nsew
rlabel metal3 19390 56060 19390 56060 0 RWL[92]
port 176 nsew
rlabel metal3 19390 56682 19390 56682 0 RWL[93]
port 177 nsew
rlabel metal3 19390 57272 19390 57272 0 RWL[94]
port 178 nsew
rlabel metal3 19390 57894 19390 57894 0 RWL[95]
port 179 nsew
rlabel metal3 19390 58484 19390 58484 0 RWL[96]
port 180 nsew
rlabel metal3 19390 59106 19390 59106 0 RWL[97]
port 181 nsew
rlabel metal3 19390 59696 19390 59696 0 RWL[98]
port 182 nsew
rlabel metal3 19390 60318 19390 60318 0 RWL[99]
port 183 nsew
rlabel metal3 19390 60908 19390 60908 0 RWL[100]
port 184 nsew
rlabel metal3 19390 61530 19390 61530 0 RWL[101]
port 185 nsew
rlabel metal3 19390 62120 19390 62120 0 RWL[102]
port 186 nsew
rlabel metal3 19390 62742 19390 62742 0 RWL[103]
port 187 nsew
rlabel metal3 19390 63332 19390 63332 0 RWL[104]
port 188 nsew
rlabel metal3 19390 63954 19390 63954 0 RWL[105]
port 189 nsew
rlabel metal3 19390 64544 19390 64544 0 RWL[106]
port 190 nsew
rlabel metal3 19390 65166 19390 65166 0 RWL[107]
port 191 nsew
rlabel metal3 19390 65756 19390 65756 0 RWL[108]
port 192 nsew
rlabel metal3 19390 66378 19390 66378 0 RWL[109]
port 193 nsew
rlabel metal3 19390 66968 19390 66968 0 RWL[110]
port 194 nsew
rlabel metal3 19390 67590 19390 67590 0 RWL[111]
port 195 nsew
rlabel metal3 19390 68180 19390 68180 0 RWL[112]
port 196 nsew
rlabel metal3 19390 68802 19390 68802 0 RWL[113]
port 197 nsew
rlabel metal3 19390 69392 19390 69392 0 RWL[114]
port 198 nsew
rlabel metal3 19390 70014 19390 70014 0 RWL[115]
port 199 nsew
rlabel metal3 19390 70604 19390 70604 0 RWL[116]
port 200 nsew
rlabel metal3 19390 71226 19390 71226 0 RWL[117]
port 201 nsew
rlabel metal3 19390 71816 19390 71816 0 RWL[118]
port 202 nsew
rlabel metal3 19390 72438 19390 72438 0 RWL[119]
port 203 nsew
rlabel metal3 19390 73028 19390 73028 0 RWL[120]
port 204 nsew
rlabel metal3 19390 73650 19390 73650 0 RWL[121]
port 205 nsew
rlabel metal3 19390 74240 19390 74240 0 RWL[122]
port 206 nsew
rlabel metal3 19390 74862 19390 74862 0 RWL[123]
port 207 nsew
rlabel metal3 19390 75452 19390 75452 0 RWL[124]
port 208 nsew
rlabel metal3 19390 76074 19390 76074 0 RWL[125]
port 209 nsew
rlabel metal3 19390 76664 19390 76664 0 RWL[126]
port 210 nsew
rlabel metal3 19390 77286 19390 77286 0 RWL[127]
port 211 nsew
rlabel metal3 44 39094 44 39094 0 LWL[64]
port 212 nsew
rlabel metal3 44 39716 44 39716 0 LWL[65]
port 213 nsew
rlabel metal3 44 40306 44 40306 0 LWL[66]
port 214 nsew
rlabel metal3 44 40928 44 40928 0 LWL[67]
port 215 nsew
rlabel metal3 44 41518 44 41518 0 LWL[68]
port 216 nsew
rlabel metal3 44 42140 44 42140 0 LWL[69]
port 217 nsew
rlabel metal3 44 42730 44 42730 0 LWL[70]
port 218 nsew
rlabel metal3 44 43352 44 43352 0 LWL[71]
port 219 nsew
rlabel metal3 44 43942 44 43942 0 LWL[72]
port 220 nsew
rlabel metal3 44 44564 44 44564 0 LWL[73]
port 221 nsew
rlabel metal3 44 45154 44 45154 0 LWL[74]
port 222 nsew
rlabel metal3 44 45776 44 45776 0 LWL[75]
port 223 nsew
rlabel metal3 44 46366 44 46366 0 LWL[76]
port 224 nsew
rlabel metal3 44 46988 44 46988 0 LWL[77]
port 225 nsew
rlabel metal3 44 47578 44 47578 0 LWL[78]
port 226 nsew
rlabel metal3 44 48200 44 48200 0 LWL[79]
port 227 nsew
rlabel metal3 44 48790 44 48790 0 LWL[80]
port 228 nsew
rlabel metal3 44 49412 44 49412 0 LWL[81]
port 229 nsew
rlabel metal3 44 50002 44 50002 0 LWL[82]
port 230 nsew
rlabel metal3 44 50624 44 50624 0 LWL[83]
port 231 nsew
rlabel metal3 44 51214 44 51214 0 LWL[84]
port 232 nsew
rlabel metal3 44 51836 44 51836 0 LWL[85]
port 233 nsew
rlabel metal3 44 52426 44 52426 0 LWL[86]
port 234 nsew
rlabel metal3 44 53048 44 53048 0 LWL[87]
port 235 nsew
rlabel metal3 44 53638 44 53638 0 LWL[88]
port 236 nsew
rlabel metal3 44 54260 44 54260 0 LWL[89]
port 237 nsew
rlabel metal3 44 54850 44 54850 0 LWL[90]
port 238 nsew
rlabel metal3 44 55472 44 55472 0 LWL[91]
port 239 nsew
rlabel metal3 44 56062 44 56062 0 LWL[92]
port 240 nsew
rlabel metal3 44 56684 44 56684 0 LWL[93]
port 241 nsew
rlabel metal3 44 57274 44 57274 0 LWL[94]
port 242 nsew
rlabel metal3 44 57896 44 57896 0 LWL[95]
port 243 nsew
rlabel metal3 44 58486 44 58486 0 LWL[96]
port 244 nsew
rlabel metal3 44 59108 44 59108 0 LWL[97]
port 245 nsew
rlabel metal3 44 59698 44 59698 0 LWL[98]
port 246 nsew
rlabel metal3 44 60320 44 60320 0 LWL[99]
port 247 nsew
rlabel metal3 44 60910 44 60910 0 LWL[100]
port 248 nsew
rlabel metal3 44 61532 44 61532 0 LWL[101]
port 249 nsew
rlabel metal3 44 62122 44 62122 0 LWL[102]
port 250 nsew
rlabel metal3 44 62744 44 62744 0 LWL[103]
port 251 nsew
rlabel metal3 44 63334 44 63334 0 LWL[104]
port 252 nsew
rlabel metal3 44 63956 44 63956 0 LWL[105]
port 253 nsew
rlabel metal3 44 64546 44 64546 0 LWL[106]
port 254 nsew
rlabel metal3 44 65168 44 65168 0 LWL[107]
port 255 nsew
rlabel metal3 44 65758 44 65758 0 LWL[108]
port 256 nsew
rlabel metal3 44 66380 44 66380 0 LWL[109]
port 257 nsew
rlabel metal3 44 66970 44 66970 0 LWL[110]
port 258 nsew
rlabel metal3 44 67592 44 67592 0 LWL[111]
port 259 nsew
rlabel metal3 44 68182 44 68182 0 LWL[112]
port 260 nsew
rlabel metal3 44 68804 44 68804 0 LWL[113]
port 261 nsew
rlabel metal3 44 69394 44 69394 0 LWL[114]
port 262 nsew
rlabel metal3 44 70016 44 70016 0 LWL[115]
port 263 nsew
rlabel metal3 44 70606 44 70606 0 LWL[116]
port 264 nsew
rlabel metal3 44 71228 44 71228 0 LWL[117]
port 265 nsew
rlabel metal3 44 71818 44 71818 0 LWL[118]
port 266 nsew
rlabel metal3 44 72440 44 72440 0 LWL[119]
port 267 nsew
rlabel metal3 44 73030 44 73030 0 LWL[120]
port 268 nsew
rlabel metal3 44 73652 44 73652 0 LWL[121]
port 269 nsew
rlabel metal3 44 74242 44 74242 0 LWL[122]
port 270 nsew
rlabel metal3 44 74864 44 74864 0 LWL[123]
port 271 nsew
rlabel metal3 44 75454 44 75454 0 LWL[124]
port 272 nsew
rlabel metal3 44 76076 44 76076 0 LWL[125]
port 273 nsew
rlabel metal3 44 76666 44 76666 0 LWL[126]
port 274 nsew
rlabel metal3 44 77288 44 77288 0 LWL[127]
port 275 nsew
<< end >>
