magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< error_s >>
rect 5257 4262 5362 4382
rect 1492 2672 1606 4262
rect 5377 3263 5482 4262
rect 6657 2672 6771 4262
<< nwell >>
rect 5170 3263 5362 5302
<< metal2 >>
rect 684 7739 775 7833
rect 933 7739 1024 7833
rect 1937 7739 2028 7833
rect 2191 7739 2282 7833
rect 2875 7014 3123 8738
rect 3650 7205 3740 8019
rect 5849 7739 5940 7833
rect 6099 7739 6189 7833
rect 7102 7739 7193 7833
rect 7356 7739 7446 7833
rect 8815 7205 8905 8019
rect 10497 7895 10744 8780
rect 9007 7640 10744 7895
rect 9007 7014 9254 7640
rect 11028 7506 11183 7991
rect 11274 7506 11429 7991
rect 12172 7506 12327 7991
rect 12418 7506 12573 7991
rect 13316 7506 13471 7991
rect 13561 7506 13717 7991
rect 14459 7506 14614 7991
rect 14705 7506 14861 7991
rect 15360 7014 15607 8738
rect 16135 7205 16226 8019
rect 3839 148 3929 242
rect 5023 148 5113 242
rect 9004 148 9095 242
rect 10187 148 10278 242
rect 16344 148 16434 242
rect 17528 148 17618 242
rect 18711 148 18802 242
<< metal3 >>
rect 32 8145 19082 8780
rect 32 7773 16226 8019
rect 5256 1563 5777 2041
rect 5256 754 5777 1390
rect 5256 0 5777 634
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_0
timestamp 1763476864
transform 1 0 3695 0 1 7896
box -44 -123 44 123
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_1
timestamp 1763476864
transform 1 0 8860 0 1 7896
box -44 -123 44 123
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_2
timestamp 1763476864
transform 1 0 16180 0 1 7896
box -44 -123 44 123
use M3_M2$$47115308_512x8m81  M3_M2$$47115308_512x8m81_0
timestamp 1763476864
transform 1 0 2979 0 1 8463
box -119 -275 119 275
use M3_M2$$47115308_512x8m81  M3_M2$$47115308_512x8m81_1
timestamp 1763476864
transform 1 0 15484 0 1 8463
box -119 -275 119 275
use M3_M2$$201412652_512x8m81  M3_M2$$201412652_512x8m81_0
timestamp 1763476864
transform 1 0 10620 0 1 8463
box -119 -275 119 275
use xpredec0_512x8m81  xpredec0_512x8m81_0
timestamp 1763476864
transform 1 0 5412 0 1 0
box -226 -1 5218 8019
use xpredec0_512x8m81  xpredec0_512x8m81_1
timestamp 1763476864
transform 1 0 247 0 1 0
box -226 -1 5218 8019
use xpredec1_512x8m81  xpredec1_512x8m81_0
timestamp 1763476864
transform 1 0 10557 0 1 0
box -1 -1 8563 7679
<< labels >>
rlabel metal3 s 15850 7917 15850 7917 4 clk
port 1 nsew
rlabel metal3 s 17852 8463 17852 8463 4 men
port 2 nsew
rlabel metal2 s 16389 195 16389 195 4 A[2]
port 3 nsew
rlabel metal2 s 3884 195 3884 195 4 A[6]
port 4 nsew
rlabel metal2 s 9049 195 9049 195 4 A[4]
port 5 nsew
rlabel metal2 s 5895 7786 5895 7786 4 xb[3]
port 6 nsew
rlabel metal2 s 14786 7945 14786 7945 4 xa[0]
port 7 nsew
rlabel metal2 s 2236 7784 2236 7784 4 xc[0]
port 8 nsew
rlabel metal2 s 1983 7784 1983 7784 4 xc[1]
port 9 nsew
rlabel metal2 s 979 7786 979 7786 4 xc[2]
port 10 nsew
rlabel metal2 s 730 7786 730 7786 4 xc[3]
port 11 nsew
rlabel metal2 s 7147 7784 7147 7784 4 xb[1]
port 12 nsew
rlabel metal2 s 6143 7786 6143 7786 4 xb[2]
port 13 nsew
rlabel metal2 s 7401 7784 7401 7784 4 xb[0]
port 14 nsew
rlabel metal2 s 14534 7945 14534 7945 4 xa[1]
port 15 nsew
rlabel metal2 s 13633 7945 13633 7945 4 xa[2]
port 16 nsew
rlabel metal2 s 13393 7945 13393 7945 4 xa[3]
port 17 nsew
rlabel metal2 s 12497 7945 12497 7945 4 xa[4]
port 18 nsew
rlabel metal2 s 12248 7945 12248 7945 4 xa[5]
port 19 nsew
rlabel metal2 s 11350 7945 11350 7945 4 xa[6]
port 20 nsew
rlabel metal2 s 11104 7945 11104 7945 4 xa[7]
port 21 nsew
rlabel metal2 s 18757 195 18757 195 4 A[0]
port 22 nsew
rlabel metal2 s 10233 195 10233 195 4 A[3]
port 23 nsew
rlabel metal2 s 5068 195 5068 195 4 A[5]
port 24 nsew
rlabel metal2 s 17573 195 17573 195 4 A[1]
port 25 nsew
<< end >>
