magic
tech gf180mcuD
magscale 1 10
timestamp 1763344618
<< metal1 >>
rect 2654 20138 4331 20232
rect 2632 16561 4157 16697
<< metal2 >>
rect 2831 25266 3510 36851
rect 2831 9963 3531 25266
rect 2831 1470 3531 9623
<< metal3 >>
rect 2337 25861 4445 26001
rect 2337 25784 3047 25861
rect 2337 25448 4445 25784
rect 2337 23893 4445 25160
rect 2337 22413 3531 23893
rect 2337 22214 4642 22413
rect 2337 20427 4445 21814
rect 3674 20424 4445 20427
rect 2337 18039 3531 18429
rect 2337 17729 4445 18039
rect 2337 16952 4445 17270
rect 2337 16570 3047 16952
rect 2337 14224 4445 16130
rect 2337 11642 4445 14024
rect 2337 11036 4445 11537
rect 2337 10605 3531 11036
rect 2337 10038 4445 10605
rect 2337 8746 4445 9668
rect 2337 7329 4445 8283
rect 2337 6510 4445 6940
rect 2337 5962 3047 6510
rect 2337 5659 4445 5962
rect 2337 5244 4445 5563
rect 2337 4783 3535 5244
rect 2337 4465 4445 4783
rect 2337 4017 4445 4263
rect 2337 3621 3037 4017
rect 2337 3374 4445 3621
rect 2337 2135 4445 2835
use M2_M14310591302080_512x8m81  M2_M14310591302080_512x8m81_0
timestamp 1763255117
transform 1 0 2648 0 1 3809
box -113 -417 113 417
use M2_M14310591302080_512x8m81  M2_M14310591302080_512x8m81_1
timestamp 1763255117
transform 1 0 2648 0 1 9199
box -113 -417 113 417
use M2_M14310591302081_512x8m81  M2_M14310591302081_512x8m81_0
timestamp 1763255117
transform 1 0 2648 0 1 16841
box -113 -330 113 330
use M2_M14310591302087_512x8m81  M2_M14310591302087_512x8m81_0
timestamp 1763255117
transform 1 0 2648 0 1 25721
box -113 -243 113 243
use M2_M14310591302092_512x8m81  M2_M14310591302092_512x8m81_0
timestamp 1763255117
transform 1 0 2648 0 1 12856
box -113 -1155 113 1155
use M2_M14310591302093_512x8m81  M2_M14310591302093_512x8m81_0
timestamp 1763255117
transform 1 0 2648 0 1 6297
box -113 -634 113 634
use M2_M14310591302093_512x8m81  M2_M14310591302093_512x8m81_1
timestamp 1763255117
transform 1 0 2648 0 1 20704
box -113 -634 113 634
use M3_M24310591302042_512x8m81  M3_M24310591302042_512x8m81_0
timestamp 1763255117
transform 1 0 3189 0 1 2483
box -330 -330 330 330
use M3_M24310591302042_512x8m81  M3_M24310591302042_512x8m81_1
timestamp 1763255117
transform 1 0 3189 0 1 18060
box -330 -330 330 330
use M3_M24310591302082_512x8m81  M3_M24310591302082_512x8m81_0
timestamp 1763255117
transform 1 0 3189 0 1 5014
box -330 -547 330 547
use M3_M24310591302083_512x8m81  M3_M24310591302083_512x8m81_0
timestamp 1763255117
transform 1 0 3189 0 1 23524
box -330 -1282 330 1632
use M3_M24310591302084_512x8m81  M3_M24310591302084_512x8m81_0
timestamp 1763255117
transform 1 0 2648 0 1 12856
box -113 -1155 113 1155
use M3_M24310591302085_512x8m81  M3_M24310591302085_512x8m81_0
timestamp 1763255117
transform 1 0 2648 0 1 16921
box -113 -330 113 330
use M3_M24310591302086_512x8m81  M3_M24310591302086_512x8m81_0
timestamp 1763255117
transform 1 0 2648 0 1 6297
box -113 -634 113 634
use M3_M24310591302086_512x8m81  M3_M24310591302086_512x8m81_1
timestamp 1763255117
transform 1 0 2648 0 1 21104
box -113 -634 113 634
use M3_M24310591302088_512x8m81  M3_M24310591302088_512x8m81_0
timestamp 1763255117
transform 1 0 3189 0 1 10795
box -330 -721 330 721
use M3_M24310591302089_512x8m81  M3_M24310591302089_512x8m81_0
timestamp 1763255117
transform 1 0 2648 0 1 3809
box -113 -417 113 417
use M3_M24310591302089_512x8m81  M3_M24310591302089_512x8m81_1
timestamp 1763255117
transform 1 0 2648 0 1 9199
box -113 -417 113 417
use M3_M24310591302090_512x8m81  M3_M24310591302090_512x8m81_0
timestamp 1763255117
transform 1 0 2648 0 1 25721
box -113 -243 113 243
use M3_M24310591302091_512x8m81  M3_M24310591302091_512x8m81_0
timestamp 1763255117
transform 1 0 3189 0 1 7800
box -330 -460 330 460
use M3_M24310591302094_512x8m81  M3_M24310591302094_512x8m81_0
timestamp 1763255117
transform 1 0 3189 0 1 15177
box -330 -938 330 938
<< end >>
