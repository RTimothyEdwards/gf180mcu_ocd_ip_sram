magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal1 >>
rect -1373 94 1373 123
rect -1373 -94 -1346 94
rect 1346 -94 1373 94
rect -1373 -123 1373 -94
<< via1 >>
rect -1346 -94 1346 94
<< metal2 >>
rect -1373 94 1373 123
rect -1373 -94 -1346 94
rect 1346 -94 1373 94
rect -1373 -122 1373 -94
<< end >>
