magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal2 >>
rect -266 172 266 198
rect -266 -172 -241 172
rect 241 -172 266 172
rect -266 -198 266 -172
<< via2 >>
rect -241 -172 241 172
<< metal3 >>
rect -266 172 266 198
rect -266 -172 -241 172
rect 241 -172 266 172
rect -266 -198 266 -172
<< end >>
