magic
tech gf180mcuD
magscale 1 10
timestamp 1763483433
<< error_s >>
rect 15574 -1957 15604 -1901
rect 15630 -1958 15660 -1957
rect 15713 -8244 15727 -8216
rect 15712 -8336 15727 -8244
<< nwell >>
rect 15513 -2147 15942 -674
rect 15513 -4026 16041 -2147
rect 15684 -7092 16041 -6739
rect 15684 -7172 16040 -7092
rect 15713 -8199 16040 -7172
rect 15713 -8316 15986 -8199
rect 15727 -8336 15986 -8316
rect 15712 -8416 15986 -8336
rect 15855 -11035 16474 -10313
rect 15876 -11036 16474 -11035
rect 15879 -14754 16477 -13599
rect 15879 -16139 16170 -15819
<< polysilicon >>
rect 16067 -10988 16123 -10969
rect 16227 -10988 16283 -10969
rect 16067 -11084 16283 -10988
rect 16067 -11181 16123 -11084
rect 16227 -11181 16283 -11084
rect 16030 -13552 16086 -13532
rect 16190 -13552 16246 -13532
rect 16030 -13644 16246 -13552
rect 16030 -13668 16086 -13644
rect 16190 -13668 16246 -13644
<< metal1 >>
rect 16572 35210 16609 35350
rect 16624 35210 16894 35350
rect -525 -240 -472 80
rect -525 -320 -275 -240
rect 16172 -3925 16353 -3213
rect 15820 -7685 16121 -7601
rect 15820 -9454 15901 -7685
rect 16357 -7970 16527 -7762
rect 15820 -9538 16522 -9454
rect 16134 -10986 16216 -10716
rect 15853 -11038 16216 -10986
rect 16440 -10996 16522 -9538
rect 15853 -13590 15904 -11038
rect 16134 -11222 16216 -11038
rect 16285 -11080 16522 -10996
rect 15977 -12861 16059 -11308
rect 15853 -13642 16062 -13590
rect 16137 -13801 16219 -12830
rect 16291 -12861 16373 -11308
rect 15981 -16021 16062 -14588
rect 16134 -16135 16225 -15948
rect 16294 -16021 16375 -14592
rect 16100 -17392 16256 -16135
<< metal2 >>
rect -528 93 -472 40214
rect 16574 38797 16661 40245
rect 16123 -599 16207 113
rect 16076 -668 16207 -599
rect 16333 -599 16417 112
rect 16574 21 16661 37818
rect 16333 -668 16422 -599
rect 16076 -795 16132 -668
rect 16366 -795 16422 -668
rect 16134 -17627 16225 -12238
<< metal3 >>
rect -631 83 -432 180
rect 15604 -1957 16729 -718
rect 15604 -1958 15630 -1957
rect 15668 -5427 16729 -4043
rect 15667 -5672 16729 -5522
rect 15667 -5918 16729 -5767
rect 15667 -6163 16729 -6012
rect 15667 -6408 16729 -6257
rect 15667 -6930 16507 -6780
rect 15667 -7172 16507 -7021
rect 15667 -7422 16507 -7272
rect 15667 -7667 16507 -7515
rect 15668 -8122 16507 -7813
rect 15668 -8900 16692 -8581
rect 15698 -11627 16382 -9720
rect 15698 -14208 16382 -11827
rect 15698 -14652 16382 -14312
rect 15645 -14814 16382 -14652
rect 15645 -15813 16382 -15245
rect 15698 -17115 16135 -16194
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_0
timestamp 1763476864
transform -1 0 99 0 1 7836
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1
timestamp 1763476864
transform -1 0 99 0 1 2988
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_2
timestamp 1763476864
transform -1 0 99 0 1 5412
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_3
timestamp 1763476864
transform -1 0 99 0 1 10260
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_4
timestamp 1763476864
transform -1 0 99 0 1 6624
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_5
timestamp 1763476864
transform -1 0 99 0 1 9048
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_6
timestamp 1763476864
transform -1 0 99 0 1 1776
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_7
timestamp 1763476864
transform -1 0 99 0 1 4200
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_8
timestamp 1763476864
transform -1 0 99 0 1 564
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_9
timestamp 1763476864
transform -1 0 99 0 1 19956
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_10
timestamp 1763476864
transform -1 0 99 0 1 23592
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_11
timestamp 1763476864
transform -1 0 99 0 1 22380
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_12
timestamp 1763476864
transform -1 0 99 0 1 24804
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_13
timestamp 1763476864
transform -1 0 99 0 1 21168
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_14
timestamp 1763476864
transform -1 0 99 0 1 12684
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_15
timestamp 1763476864
transform -1 0 99 0 1 17532
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_16
timestamp 1763476864
transform -1 0 99 0 1 15108
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_17
timestamp 1763476864
transform -1 0 99 0 1 16320
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_18
timestamp 1763476864
transform -1 0 99 0 1 18744
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_19
timestamp 1763476864
transform -1 0 99 0 1 13896
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_20
timestamp 1763476864
transform -1 0 99 0 1 28440
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_21
timestamp 1763476864
transform -1 0 99 0 1 30864
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_22
timestamp 1763476864
transform -1 0 99 0 1 33288
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_23
timestamp 1763476864
transform -1 0 99 0 1 38136
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_24
timestamp 1763476864
transform -1 0 99 0 1 35712
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_25
timestamp 1763476864
transform -1 0 99 0 1 27228
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_26
timestamp 1763476864
transform -1 0 99 0 1 29652
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_27
timestamp 1763476864
transform -1 0 99 0 1 32076
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_28
timestamp 1763476864
transform -1 0 99 0 1 36924
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_29
timestamp 1763476864
transform -1 0 99 0 1 34500
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_30
timestamp 1763476864
transform -1 0 99 0 1 26016
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_31
timestamp 1763476864
transform -1 0 99 0 1 11472
box 62 103 538 1445
use 018SRAM_cell1_512x8m81  018SRAM_cell1_512x8m81_0
timestamp 1763476864
transform -1 0 99 0 1 0
box 62 89 538 797
use 018SRAM_cell1_512x8m81  018SRAM_cell1_512x8m81_1
timestamp 1763476864
transform -1 0 99 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_0
timestamp 1763476864
transform -1 0 11822 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_1
timestamp 1763476864
transform -1 0 11386 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_2
timestamp 1763476864
transform -1 0 10950 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_3
timestamp 1763476864
transform -1 0 10514 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_4
timestamp 1763476864
transform -1 0 9642 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_5
timestamp 1763476864
transform -1 0 10078 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_6
timestamp 1763476864
transform -1 0 9206 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_7
timestamp 1763476864
transform -1 0 8770 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_8
timestamp 1763476864
transform -1 0 12678 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_9
timestamp 1763476864
transform -1 0 13114 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_10
timestamp 1763476864
transform -1 0 13986 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_11
timestamp 1763476864
transform -1 0 13550 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_12
timestamp 1763476864
transform -1 0 14422 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_13
timestamp 1763476864
transform -1 0 14858 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_14
timestamp 1763476864
transform -1 0 15294 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_15
timestamp 1763476864
transform -1 0 15730 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_16
timestamp 1763476864
transform -1 0 5298 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_17
timestamp 1763476864
transform -1 0 6170 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_18
timestamp 1763476864
transform -1 0 5734 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_19
timestamp 1763476864
transform -1 0 6606 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_20
timestamp 1763476864
transform -1 0 7042 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_21
timestamp 1763476864
transform -1 0 7478 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_22
timestamp 1763476864
transform -1 0 7914 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_23
timestamp 1763476864
transform -1 0 4006 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_24
timestamp 1763476864
transform -1 0 3570 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_25
timestamp 1763476864
transform -1 0 3134 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_26
timestamp 1763476864
transform -1 0 2698 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_27
timestamp 1763476864
transform -1 0 1826 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_28
timestamp 1763476864
transform -1 0 2262 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_29
timestamp 1763476864
transform -1 0 1390 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_30
timestamp 1763476864
transform -1 0 954 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_31
timestamp 1763476864
transform -1 0 4862 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_32
timestamp 1763476864
transform -1 0 2698 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_33
timestamp 1763476864
transform -1 0 1826 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_34
timestamp 1763476864
transform -1 0 2262 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_35
timestamp 1763476864
transform -1 0 1390 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_36
timestamp 1763476864
transform -1 0 954 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_37
timestamp 1763476864
transform -1 0 3570 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_38
timestamp 1763476864
transform -1 0 3134 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_39
timestamp 1763476864
transform -1 0 7478 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_40
timestamp 1763476864
transform -1 0 4862 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_41
timestamp 1763476864
transform -1 0 7914 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_42
timestamp 1763476864
transform -1 0 5298 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_43
timestamp 1763476864
transform -1 0 6170 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_44
timestamp 1763476864
transform -1 0 5734 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_45
timestamp 1763476864
transform -1 0 6606 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_46
timestamp 1763476864
transform -1 0 7042 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_47
timestamp 1763476864
transform -1 0 4006 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_48
timestamp 1763476864
transform -1 0 9642 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_49
timestamp 1763476864
transform -1 0 11386 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_50
timestamp 1763476864
transform -1 0 8770 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_51
timestamp 1763476864
transform -1 0 9206 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_52
timestamp 1763476864
transform -1 0 11822 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_53
timestamp 1763476864
transform -1 0 10078 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_54
timestamp 1763476864
transform -1 0 10514 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_55
timestamp 1763476864
transform -1 0 10950 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_56
timestamp 1763476864
transform -1 0 13550 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_57
timestamp 1763476864
transform -1 0 13114 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_59
timestamp 1763476864
transform -1 0 14422 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_60
timestamp 1763476864
transform -1 0 15294 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_61
timestamp 1763476864
transform -1 0 13986 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_62
timestamp 1763476864
transform -1 0 15730 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_63
timestamp 1763476864
transform -1 0 12678 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_64
timestamp 1763476864
transform -1 0 14858 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_0
timestamp 1763476864
transform 1 0 15986 0 -1 5100
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_1
timestamp 1763476864
transform 1 0 15986 0 -1 6312
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_2
timestamp 1763476864
transform 1 0 15986 0 -1 3888
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_3
timestamp 1763476864
transform 1 0 15986 0 -1 2676
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_4
timestamp 1763476864
transform 1 0 15986 0 -1 7524
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_5
timestamp 1763476864
transform 1 0 15986 0 -1 12372
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_6
timestamp 1763476864
transform 1 0 15986 0 -1 11160
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_7
timestamp 1763476864
transform 1 0 15986 0 -1 9948
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_8
timestamp 1763476864
transform 1 0 15986 0 -1 8736
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_9
timestamp 1763476864
transform 1 0 15986 0 -1 1464
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_10
timestamp 1763476864
transform 1 0 15986 0 1 3636
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_11
timestamp 1763476864
transform 1 0 15986 0 1 4848
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_12
timestamp 1763476864
transform 1 0 15986 0 1 7272
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_13
timestamp 1763476864
transform 1 0 15986 0 1 9696
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_14
timestamp 1763476864
transform 1 0 15986 0 1 2424
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_15
timestamp 1763476864
transform 1 0 15986 0 1 6060
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_16
timestamp 1763476864
transform 1 0 15986 0 1 8484
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_17
timestamp 1763476864
transform 1 0 15986 0 1 10908
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_18
timestamp 1763476864
transform 1 0 15986 0 1 1212
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_19
timestamp 1763476864
transform 1 0 15986 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_20
timestamp 1763476864
transform 1 0 15986 0 -1 25704
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_21
timestamp 1763476864
transform 1 0 15986 0 -1 20856
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_22
timestamp 1763476864
transform 1 0 15986 0 -1 24492
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_23
timestamp 1763476864
transform 1 0 15986 0 -1 23280
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_24
timestamp 1763476864
transform 1 0 15986 0 -1 22068
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_25
timestamp 1763476864
transform 1 0 15986 0 -1 16008
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_26
timestamp 1763476864
transform 1 0 15986 0 -1 13584
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_27
timestamp 1763476864
transform 1 0 15986 0 -1 14796
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_28
timestamp 1763476864
transform 1 0 15986 0 -1 19644
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_29
timestamp 1763476864
transform 1 0 15986 0 -1 18432
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_30
timestamp 1763476864
transform 1 0 15986 0 -1 17220
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_31
timestamp 1763476864
transform 1 0 15986 0 1 24240
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_32
timestamp 1763476864
transform 1 0 15986 0 1 20604
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_33
timestamp 1763476864
transform 1 0 15986 0 1 14544
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_34
timestamp 1763476864
transform 1 0 15986 0 1 16968
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_35
timestamp 1763476864
transform 1 0 15986 0 1 19392
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_36
timestamp 1763476864
transform 1 0 15986 0 1 21816
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_37
timestamp 1763476864
transform 1 0 15986 0 1 23028
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_38
timestamp 1763476864
transform 1 0 15986 0 1 13332
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_39
timestamp 1763476864
transform 1 0 15986 0 1 15756
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_40
timestamp 1763476864
transform 1 0 15986 0 1 18180
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_41
timestamp 1763476864
transform 1 0 15986 0 1 25452
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_42
timestamp 1763476864
transform 1 0 15986 0 -1 37824
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_43
timestamp 1763476864
transform 1 0 15986 0 -1 35400
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_44
timestamp 1763476864
transform 1 0 15986 0 -1 32976
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_45
timestamp 1763476864
transform 1 0 15986 0 -1 29340
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_46
timestamp 1763476864
transform 1 0 15986 0 -1 28128
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_47
timestamp 1763476864
transform 1 0 15986 0 -1 39036
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_48
timestamp 1763476864
transform 1 0 15986 0 -1 36612
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_49
timestamp 1763476864
transform 1 0 15986 0 -1 34188
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_50
timestamp 1763476864
transform 1 0 15986 0 -1 31764
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_51
timestamp 1763476864
transform 1 0 15986 0 -1 30552
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_52
timestamp 1763476864
transform 1 0 15986 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_53
timestamp 1763476864
transform 1 0 15986 0 1 36360
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_54
timestamp 1763476864
transform 1 0 15986 0 1 26664
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_55
timestamp 1763476864
transform 1 0 15986 0 1 31512
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_56
timestamp 1763476864
transform 1 0 15986 0 1 37572
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_57
timestamp 1763476864
transform 1 0 15986 0 1 33936
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_58
timestamp 1763476864
transform 1 0 15986 0 1 29088
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_59
timestamp 1763476864
transform 1 0 15986 0 1 38784
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_60
timestamp 1763476864
transform 1 0 15986 0 1 30300
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_61
timestamp 1763476864
transform 1 0 15986 0 1 35148
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_62
timestamp 1763476864
transform 1 0 15986 0 1 27876
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_63
timestamp 1763476864
transform 1 0 15986 0 1 32724
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_64
timestamp 1763476864
transform 1 0 15986 0 -1 26916
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_65
timestamp 1763476864
transform 1 0 15986 0 1 12120
box 62 89 538 797
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_0
timestamp 1763476864
transform -1 0 12251 0 1 0
box 91 55 511 797
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_1
timestamp 1763476864
transform -1 0 4435 0 1 0
box 91 55 511 797
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_2
timestamp 1763476864
transform -1 0 527 0 1 0
box 91 55 511 797
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_3
timestamp 1763476864
transform -1 0 4435 0 -1 40248
box 91 55 511 797
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_4
timestamp 1763476864
transform -1 0 12251 0 -1 40248
box 91 55 511 797
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_5
timestamp 1763476864
transform 1 0 15557 0 -1 40248
box 91 55 511 797
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_6
timestamp 1763476864
transform -1 0 8343 0 1 0
box 91 55 511 797
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_7
timestamp 1763476864
transform -1 0 8343 0 -1 40248
box 91 55 511 797
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_0
timestamp 1763476864
transform 1 0 15557 0 1 0
box 91 55 511 797
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_54
timestamp 1763476864
transform -1 0 527 0 -1 40248
box 91 55 511 797
use M1_NWELL$$44998700_512x8m81  M1_NWELL$$44998700_512x8m81_0
timestamp 1763476864
transform 1 0 16322 0 1 -15979
box -154 -159 154 159
use M1_NWELL$$44998700_512x8m81  M1_NWELL$$44998700_512x8m81_1
timestamp 1763476864
transform 1 0 15941 0 1 -15979
box -154 -159 154 159
use M1_NWELL$$46277676_512x8m81  M1_NWELL$$46277676_512x8m81_0
timestamp 1763476864
transform 1 0 16135 0 1 -10155
box -265 -159 265 159
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_0
timestamp 1763476864
transform 1 0 16620 0 -1 4974
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_1
timestamp 1763476864
transform 1 0 16620 0 -1 3762
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_2
timestamp 1763476864
transform 1 0 16620 0 -1 1338
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_3
timestamp 1763476864
transform 1 0 16620 0 -1 126
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_4
timestamp 1763476864
transform 1 0 16620 0 -1 11034
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_5
timestamp 1763476864
transform 1 0 16620 0 -1 8610
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_6
timestamp 1763476864
transform 1 0 16620 0 -1 6186
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_7
timestamp 1763476864
transform 1 0 16620 0 -1 9822
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_8
timestamp 1763476864
transform 1 0 16620 0 -1 7398
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_9
timestamp 1763476864
transform 1 0 16620 0 -1 2550
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_10
timestamp 1763476864
transform 1 0 16620 0 -1 14670
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_11
timestamp 1763476864
transform 1 0 16620 0 -1 25578
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_12
timestamp 1763476864
transform 1 0 16620 0 -1 24366
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_13
timestamp 1763476864
transform 1 0 16620 0 -1 23154
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_14
timestamp 1763476864
transform 1 0 16620 0 -1 21942
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_15
timestamp 1763476864
transform 1 0 16620 0 -1 20730
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_16
timestamp 1763476864
transform 1 0 16620 0 -1 18306
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_17
timestamp 1763476864
transform 1 0 16620 0 -1 15882
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_18
timestamp 1763476864
transform 1 0 16620 0 -1 13458
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_19
timestamp 1763476864
transform 1 0 16620 0 -1 19518
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_20
timestamp 1763476864
transform 1 0 16620 0 -1 17094
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_21
timestamp 1763476864
transform 1 0 16620 0 -1 37698
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_22
timestamp 1763476864
transform 1 0 16620 0 -1 36486
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_23
timestamp 1763476864
transform 1 0 16620 0 -1 35274
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_24
timestamp 1763476864
transform 1 0 16620 0 -1 34062
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_25
timestamp 1763476864
transform 1 0 16620 0 -1 32850
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_26
timestamp 1763476864
transform 1 0 16620 0 -1 31638
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_27
timestamp 1763476864
transform 1 0 16620 0 -1 30426
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_28
timestamp 1763476864
transform 1 0 16620 0 -1 29214
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_29
timestamp 1763476864
transform 1 0 16620 0 -1 28002
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_30
timestamp 1763476864
transform 1 0 16620 0 -1 26790
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_31
timestamp 1763476864
transform 1 0 16620 0 -1 38910
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_32
timestamp 1763476864
transform 1 0 16620 0 -1 40122
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_33
timestamp 1763476864
transform 1 0 16620 0 -1 12246
box -96 -124 67 124
use M1_POLY2$$46559276_512x8m81_0  M1_POLY2$$46559276_512x8m81_0_0
timestamp 1763476864
transform -1 0 15966 0 1 -13600
box -123 -48 123 48
use M1_POLY2$$46559276_512x8m81_0  M1_POLY2$$46559276_512x8m81_0_1
timestamp 1763476864
transform 1 0 16375 0 1 -11038
box -123 -48 123 48
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_0
timestamp 1763476864
transform 1 0 -499 0 1 128
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_1
timestamp 1763476864
transform 1 0 -499 0 1 1340
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_2
timestamp 1763476864
transform 1 0 -499 0 1 2552
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_3
timestamp 1763476864
transform 1 0 -499 0 1 4976
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_4
timestamp 1763476864
transform 1 0 -499 0 1 3764
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_5
timestamp 1763476864
transform 1 0 -499 0 1 9824
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_6
timestamp 1763476864
transform 1 0 -499 0 1 8612
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_7
timestamp 1763476864
transform 1 0 -499 0 1 11036
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_8
timestamp 1763476864
transform 1 0 -499 0 1 12248
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_9
timestamp 1763476864
transform 1 0 -499 0 1 7400
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_10
timestamp 1763476864
transform 1 0 -499 0 1 6188
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_11
timestamp 1763476864
transform 1 0 -499 0 1 14672
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_12
timestamp 1763476864
transform 1 0 -499 0 1 13460
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_13
timestamp 1763476864
transform 1 0 -499 0 1 15884
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_14
timestamp 1763476864
transform 1 0 -499 0 1 17096
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_15
timestamp 1763476864
transform 1 0 -499 0 1 19520
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_16
timestamp 1763476864
transform 1 0 -499 0 1 18308
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_17
timestamp 1763476864
transform 1 0 -499 0 1 20732
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_18
timestamp 1763476864
transform 1 0 -499 0 1 21944
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_19
timestamp 1763476864
transform 1 0 -499 0 1 24368
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_20
timestamp 1763476864
transform 1 0 -499 0 1 23156
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_21
timestamp 1763476864
transform 1 0 -499 0 1 25580
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_22
timestamp 1763476864
transform 1 0 -499 0 1 26792
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_23
timestamp 1763476864
transform 1 0 -499 0 1 29216
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_24
timestamp 1763476864
transform 1 0 -499 0 1 28004
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_25
timestamp 1763476864
transform 1 0 -499 0 1 30428
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_26
timestamp 1763476864
transform 1 0 -499 0 1 31640
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_27
timestamp 1763476864
transform 1 0 -499 0 1 34064
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_28
timestamp 1763476864
transform 1 0 -499 0 1 32852
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_29
timestamp 1763476864
transform 1 0 -499 0 1 35276
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_30
timestamp 1763476864
transform 1 0 -499 0 1 36488
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_31
timestamp 1763476864
transform 1 0 -499 0 1 38912
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_32
timestamp 1763476864
transform 1 0 -499 0 1 37700
box -36 -126 60 122
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_33
timestamp 1763476864
transform 1 0 -499 0 1 40124
box -36 -126 60 122
use M1_PSUB$$46274604_512x8m81  M1_PSUB$$46274604_512x8m81_0
timestamp 1763476864
transform 1 0 16174 0 1 -11551
box -166 -58 166 58
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1763476864
transform 1 0 16618 0 -1 11034
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_1
timestamp 1763476864
transform 1 0 16618 0 -1 8610
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_2
timestamp 1763476864
transform 1 0 16618 0 -1 6185
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_3
timestamp 1763476864
transform 1 0 16618 0 -1 3761
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_4
timestamp 1763476864
transform 1 0 16618 0 -1 1339
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_5
timestamp 1763476864
transform 1 0 16618 0 -1 7398
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_6
timestamp 1763476864
transform 1 0 16618 0 -1 2550
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_7
timestamp 1763476864
transform 1 0 16618 0 -1 127
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_8
timestamp 1763476864
transform 1 0 16618 0 -1 9825
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_9
timestamp 1763476864
transform 1 0 16618 0 -1 4974
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_10
timestamp 1763476864
transform 1 0 16618 0 -1 21942
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_11
timestamp 1763476864
transform 1 0 16618 0 -1 20730
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_12
timestamp 1763476864
transform 1 0 16618 0 -1 18306
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_13
timestamp 1763476864
transform 1 0 16618 0 -1 15882
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_14
timestamp 1763476864
transform 1 0 16618 0 -1 13458
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_15
timestamp 1763476864
transform 1 0 16618 0 -1 17097
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_16
timestamp 1763476864
transform 1 0 16618 0 -1 19518
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_17
timestamp 1763476864
transform 1 0 16618 0 -1 25578
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_18
timestamp 1763476864
transform 1 0 16618 0 -1 14673
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_19
timestamp 1763476864
transform 1 0 16618 0 -1 24366
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_20
timestamp 1763476864
transform 1 0 16618 0 -1 23154
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_21
timestamp 1763476864
transform 1 0 16618 0 -1 37698
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_22
timestamp 1763476864
transform 1 0 16618 0 -1 36486
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_23
timestamp 1763476864
transform 1 0 16618 0 -1 35274
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_24
timestamp 1763476864
transform 1 0 16618 0 -1 34062
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_25
timestamp 1763476864
transform 1 0 16618 0 -1 32850
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_26
timestamp 1763476864
transform 1 0 16618 0 -1 31638
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_27
timestamp 1763476864
transform 1 0 16618 0 -1 30426
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_28
timestamp 1763476864
transform 1 0 16618 0 -1 29214
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_29
timestamp 1763476864
transform 1 0 16618 0 -1 28002
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_30
timestamp 1763476864
transform 1 0 16618 0 -1 26790
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_31
timestamp 1763476864
transform 1 0 16618 0 -1 40122
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_32
timestamp 1763476864
transform 1 0 16618 0 -1 38910
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_33
timestamp 1763476864
transform 1 0 16618 0 -1 12249
box -43 -122 43 122
use M2_M1$$47117356_512x8m81  M2_M1$$47117356_512x8m81_0
timestamp 1763476864
transform 1 0 16179 0 1 -14108
box -45 -1874 45 1874
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_0
timestamp 1763476864
transform 1 0 -499 0 1 1340
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_1
timestamp 1763476864
transform 1 0 -499 0 1 2552
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_2
timestamp 1763476864
transform 1 0 -499 0 1 3764
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_3
timestamp 1763476864
transform 1 0 -499 0 1 4976
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_4
timestamp 1763476864
transform 1 0 -499 0 1 6188
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_5
timestamp 1763476864
transform 1 0 -499 0 1 7400
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_6
timestamp 1763476864
transform 1 0 -499 0 1 8612
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_7
timestamp 1763476864
transform 1 0 -499 0 1 9824
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_8
timestamp 1763476864
transform 1 0 -499 0 1 11036
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_9
timestamp 1763476864
transform 1 0 -499 0 1 12248
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_10
timestamp 1763476864
transform 1 0 -499 0 1 25580
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_11
timestamp 1763476864
transform 1 0 -499 0 1 24368
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_12
timestamp 1763476864
transform 1 0 -499 0 1 23156
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_13
timestamp 1763476864
transform 1 0 -499 0 1 21944
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_14
timestamp 1763476864
transform 1 0 -499 0 1 20732
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_15
timestamp 1763476864
transform 1 0 -499 0 1 19520
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_16
timestamp 1763476864
transform 1 0 -499 0 1 18308
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_17
timestamp 1763476864
transform 1 0 -499 0 1 17096
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_18
timestamp 1763476864
transform 1 0 -499 0 1 13460
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_19
timestamp 1763476864
transform 1 0 -499 0 1 14672
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_20
timestamp 1763476864
transform 1 0 -502 0 1 15884
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_21
timestamp 1763476864
transform 1 0 -499 0 1 38911
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_22
timestamp 1763476864
transform 1 0 -499 0 1 37700
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_23
timestamp 1763476864
transform 1 0 -499 0 1 36488
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_24
timestamp 1763476864
transform 1 0 -499 0 1 35276
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_25
timestamp 1763476864
transform 1 0 -499 0 1 34063
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_26
timestamp 1763476864
transform 1 0 -499 0 1 32852
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_27
timestamp 1763476864
transform 1 0 -499 0 1 31640
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_28
timestamp 1763476864
transform 1 0 -499 0 1 30428
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_29
timestamp 1763476864
transform 1 0 -499 0 1 29216
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_30
timestamp 1763476864
transform 1 0 -499 0 1 28004
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_31
timestamp 1763476864
transform 1 0 -499 0 1 26792
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_32
timestamp 1763476864
transform 1 0 -499 0 1 40081
box -34 -99 34 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_0
timestamp 1763476864
transform 0 -1 -532 1 0 128
box -35 -99 35 99
use nmos_5p04310591302096_512x8m81  nmos_5p04310591302096_512x8m81_0
timestamp 1763476864
transform 1 0 16058 0 1 -13502
box -116 -44 276 837
use nmos_5p04310591302098_512x8m81  nmos_5p04310591302098_512x8m81_0
timestamp 1763476864
transform 1 0 16095 0 1 -11342
box -116 -44 276 172
use pmos_5p04310591302095_512x8m81  pmos_5p04310591302095_512x8m81_0
timestamp 1763476864
transform 1 0 16095 0 1 -10936
box -202 -86 362 413
use pmos_5p04310591302097_512x8m81  pmos_5p04310591302097_512x8m81_0
timestamp 1763476864
transform 1 0 16058 0 -1 -13698
box -202 -86 362 1079
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_0
timestamp 1763476864
transform 1 0 16298 0 1 -12832
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_1
timestamp 1763476864
transform 1 0 16299 0 1 -10749
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_2
timestamp 1763476864
transform 1 0 16301 0 1 -15787
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_3
timestamp 1763476864
transform 1 0 15992 0 1 -15507
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_4
timestamp 1763476864
transform 1 0 15989 0 1 -12456
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_5
timestamp 1763476864
transform 1 0 15989 0 1 -13256
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_6
timestamp 1763476864
transform 1 0 15985 0 1 -10749
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_7
timestamp 1763476864
transform 1 0 16301 0 1 -15507
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_8
timestamp 1763476864
transform 1 0 15989 0 1 -12832
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_9
timestamp 1763476864
transform 1 0 15992 0 1 -15787
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_10
timestamp 1763476864
transform 1 0 16298 0 1 -12456
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_11
timestamp 1763476864
transform 1 0 16298 0 1 -13256
box -9 0 73 215
use via1_2_x2_R90_512x8m81_0  via1_2_x2_R90_512x8m81_0_0
timestamp 1763476864
transform 0 -1 16230 1 0 -10189
box -9 0 73 215
use via1_2_x2_R270_512x8m81_0  via1_2_x2_R270_512x8m81_0_0
timestamp 1763476864
transform 0 1 15995 -1 0 -7771
box -9 0 75 215
use ypass_gate_512x8m81_0  ypass_gate_512x8m81_0_0
timestamp 1763482574
transform -1 0 16476 0 1 -9333
box -155 371 651 8659
<< end >>
