magic
tech gf180mcuD
magscale 1 10
timestamp 1763485967
<< nwell >>
rect -32 10266 602 11861
rect -7 9396 602 10266
rect -5 8409 602 9396
rect -5 4480 633 4880
rect -13 4475 633 4480
rect -130 4019 633 4475
<< pmos >>
rect 172 10921 228 11239
rect 332 10921 388 11239
rect 172 10416 228 10733
rect 332 10416 388 10733
rect 169 4108 225 4247
rect 376 4108 432 4247
<< ndiff >>
rect 54 3843 80 3915
rect 489 3843 505 3915
<< pdiff >>
rect 54 11195 172 11239
rect 54 11149 97 11195
rect 143 11149 172 11195
rect 54 11013 172 11149
rect 54 10967 97 11013
rect 143 10967 172 11013
rect 54 10921 172 10967
rect 228 11195 332 11239
rect 228 11149 257 11195
rect 303 11149 332 11195
rect 228 11013 332 11149
rect 228 10967 257 11013
rect 303 10967 332 11013
rect 228 10921 332 10967
rect 388 11195 505 11239
rect 388 11149 419 11195
rect 465 11149 505 11195
rect 388 11013 505 11149
rect 388 10967 419 11013
rect 465 10967 505 11013
rect 388 10921 505 10967
rect 54 10690 172 10733
rect 54 10644 97 10690
rect 143 10644 172 10690
rect 54 10508 172 10644
rect 54 10462 97 10508
rect 143 10462 172 10508
rect 54 10416 172 10462
rect 228 10690 332 10733
rect 228 10644 257 10690
rect 303 10644 332 10690
rect 228 10508 332 10644
rect 228 10462 257 10508
rect 303 10462 332 10508
rect 228 10416 332 10462
rect 388 10690 505 10733
rect 388 10644 419 10690
rect 465 10644 505 10690
rect 388 10508 505 10644
rect 388 10462 419 10508
rect 465 10462 505 10508
rect 388 10416 505 10462
rect 36 4202 169 4247
rect 36 4155 78 4202
rect 124 4155 169 4202
rect 36 4108 169 4155
rect 225 4201 376 4247
rect 225 4155 280 4201
rect 326 4155 376 4201
rect 225 4108 376 4155
rect 432 4201 547 4247
rect 432 4155 482 4201
rect 528 4155 547 4201
rect 432 4108 547 4155
<< pdiffc >>
rect 97 11149 143 11195
rect 97 10967 143 11013
rect 257 11149 303 11195
rect 257 10967 303 11013
rect 419 11149 465 11195
rect 419 10967 465 11013
rect 97 10644 143 10690
rect 97 10462 143 10508
rect 257 10644 303 10690
rect 257 10462 303 10508
rect 419 10644 465 10690
rect 419 10462 465 10508
rect 78 4155 124 4202
rect 280 4155 326 4201
rect 482 4155 528 4201
<< nsubdiff >>
rect 119 11552 516 11712
<< polysilicon >>
rect 172 11239 228 11436
rect 332 11239 388 11436
rect 172 10733 228 10921
rect 332 10733 388 10921
rect 172 10352 228 10416
rect 332 10352 388 10416
rect 172 10268 388 10352
rect 172 10267 304 10268
rect 248 10118 304 10267
rect 250 8479 306 8553
rect 250 8400 315 8479
rect 250 6868 306 7515
rect 250 5995 306 6148
rect 250 5645 306 5852
rect 169 4386 432 4485
rect 169 4247 225 4386
rect 376 4247 432 4386
rect 169 4083 225 4108
rect 169 4010 228 4083
rect 376 4072 432 4108
rect 172 3950 228 4010
rect 340 4010 432 4072
rect 340 3950 396 4010
rect 172 3781 228 3810
rect 340 3781 396 3810
<< metal1 >>
rect 50 11562 510 11717
rect 77 11434 480 11562
rect 77 11195 159 11434
rect 77 11149 97 11195
rect 143 11149 159 11195
rect 77 11013 159 11149
rect 77 10967 97 11013
rect 143 10967 159 11013
rect 77 10690 159 10967
rect 222 11195 337 11382
rect 222 11149 257 11195
rect 303 11149 337 11195
rect 222 11013 337 11149
rect 222 10967 257 11013
rect 303 10967 337 11013
rect 222 10930 337 10967
rect 402 11195 480 11434
rect 402 11149 419 11195
rect 465 11149 480 11195
rect 402 11013 480 11149
rect 402 10967 419 11013
rect 465 10967 480 11013
rect 77 10644 97 10690
rect 143 10644 159 10690
rect 77 10508 159 10644
rect 77 10462 97 10508
rect 143 10462 159 10508
rect 77 10425 159 10462
rect 222 10690 337 10879
rect 222 10644 257 10690
rect 303 10644 337 10690
rect 222 10508 337 10644
rect 222 10462 257 10508
rect 303 10462 337 10508
rect 222 10425 337 10462
rect 402 10690 480 10967
rect 402 10644 419 10690
rect 465 10644 480 10690
rect 402 10508 480 10644
rect 402 10462 419 10508
rect 465 10462 480 10508
rect 402 10425 480 10462
rect 88 9710 219 9890
rect 333 9710 463 9890
rect 88 9066 182 9240
rect 138 8750 182 9066
rect 119 8673 182 8750
rect 381 9075 463 9240
rect 119 7560 189 8673
rect 239 8296 315 8480
rect 381 7478 465 9075
rect 45 7381 465 7478
rect 43 7103 506 7237
rect 123 6938 466 7035
rect 123 6191 188 6938
rect 380 6233 433 6816
rect 123 5665 180 6191
rect 247 5939 328 6074
rect 247 5773 328 5884
rect 123 4971 181 5665
rect 378 4818 433 6233
rect 54 4202 131 4693
rect 199 4396 329 4493
rect 54 4155 78 4202
rect 124 4155 131 4202
rect 54 4117 131 4155
rect 245 4201 328 4317
rect 245 4155 280 4201
rect 326 4155 328 4201
rect 53 3742 157 3971
rect 245 3851 328 4155
rect 466 4201 537 4693
rect 466 4155 482 4201
rect 528 4155 537 4201
rect 466 4117 537 4155
rect 415 3742 505 3971
rect 53 3470 505 3742
<< metal2 >>
rect 88 11314 144 11715
rect 216 11435 344 11717
rect 245 11434 344 11435
rect 88 11258 327 11314
rect 88 9109 144 11258
rect 421 10808 477 11715
rect 285 10752 477 10808
rect 26 7394 129 7464
rect 26 3470 82 7394
rect 248 7338 304 8406
rect 138 7282 304 7338
rect 138 5865 194 7282
rect 421 6929 477 10752
rect 381 6074 444 6848
rect 260 5977 444 6074
rect 138 5838 245 5865
rect 138 5782 312 5838
rect 138 5754 245 5782
rect 138 4317 194 5754
rect 381 5094 444 5977
rect 250 4997 444 5094
rect 250 4386 306 4997
rect 138 4138 326 4317
rect 138 4137 290 4138
rect 172 3520 272 3749
<< metal3 >>
rect -65 10338 525 11716
rect -41 7007 525 8407
rect -41 6761 525 6901
rect -41 6519 525 6659
rect -41 6278 525 6418
rect -41 6036 525 6176
rect -41 5504 525 5644
rect -41 5262 525 5402
rect -41 5020 525 5160
rect -41 4778 525 4918
rect -41 4190 525 4632
rect -41 3519 525 3974
use M1_NWELL05_512x8m81  M1_NWELL05_512x8m81_0
timestamp 1763476864
transform 1 0 285 0 1 11632
box -265 -159 265 159
use M1_NWELL09_512x8m81  M1_NWELL09_512x8m81_1
timestamp 1763476864
transform 1 0 287 0 1 4633
box -320 -159 320 159
use M1_POLY24310591302030_512x8m81  M1_POLY24310591302030_512x8m81_0
timestamp 1763476864
transform 1 0 272 0 1 10310
box -95 -36 95 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1763476864
transform 1 0 253 0 1 4443
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1763476864
transform 1 0 290 0 1 5810
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_2
timestamp 1763476864
transform 1 0 281 0 1 6037
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_6
timestamp 1763476864
transform 1 0 276 0 1 8442
box -36 -36 36 36
use M1_PSUB$$45111340_512x8m81  M1_PSUB$$45111340_512x8m81_0
timestamp 1763476864
transform 1 0 150 0 1 7168
box -56 -58 56 58
use M1_PSUB$$47122476_512x8m81  M1_PSUB$$47122476_512x8m81_0
timestamp 1763476864
transform 1 0 277 0 1 3544
box -223 -58 254 57
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_0
timestamp 1763476864
transform 1 0 287 0 1 4227
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_2
timestamp 1763476864
transform 1 0 122 0 1 9800
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_3
timestamp 1763476864
transform 1 0 122 0 1 9171
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_4
timestamp 1763476864
transform 1 0 281 0 1 11285
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_5
timestamp 1763476864
transform 1 0 276 0 1 8389
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_6
timestamp 1763476864
transform 1 0 430 0 1 9800
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_7
timestamp 1763476864
transform 1 0 281 0 1 10780
box -34 -63 34 63
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_0
timestamp 1763476864
transform 1 0 285 0 1 4442
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_1
timestamp 1763476864
transform 1 0 280 0 1 5810
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_5
timestamp 1763476864
transform 0 -1 120 1 0 7429
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_6
timestamp 1763476864
transform 1 0 324 0 1 7162
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_9
timestamp 1763476864
transform 1 0 436 0 1 6984
box -35 -56 35 55
use M3_M2431059130201_512x8m81  M3_M2431059130201_512x8m81_1
timestamp 1763476864
transform 1 0 324 0 1 7157
box -35 -63 35 63
use nmos_1p2$$47119404_512x8m81  nmos_1p2$$47119404_512x8m81_1
timestamp 1763476864
transform 1 0 264 0 -1 6826
box -102 -44 130 679
use nmos_1p2$$47119404_512x8m81  nmos_1p2$$47119404_512x8m81_3
timestamp 1763476864
transform 1 0 264 0 -1 8190
box -102 -44 130 679
use nmos_5p0431059130202_512x8m81  nmos_5p0431059130202_512x8m81_0
timestamp 1763476864
transform 1 0 204 0 1 3853
box -124 -44 285 98
use pmos_1p2$$46889004_512x8m81  pmos_1p2$$46889004_512x8m81_1
timestamp 1763476864
transform 1 0 264 0 -1 5601
box -188 -86 216 721
use pmos_5p0431059130201_512x8m81  pmos_5p0431059130201_512x8m81_0
timestamp 1763476864
transform 1 0 248 0 -1 10077
box -174 -86 230 721
use pmos_5p0431059130201_512x8m81  pmos_5p0431059130201_512x8m81_1
timestamp 1763476864
transform 1 0 250 0 -1 9231
box -174 -86 230 721
use via1_2_512x8m81  via1_2_512x8m81_0
timestamp 1763476864
transform 1 0 174 0 1 3559
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_0
timestamp 1763476864
transform -1 0 328 0 -1 6067
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_2
timestamp 1763476864
transform 0 -1 343 1 0 11435
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_3
timestamp 1763476864
transform 0 -1 343 1 0 11621
box 0 0 65 89
use via2_R90_512x8m81  via2_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 333 1 0 11435
box 0 0 65 89
use via2_R90_512x8m81  via2_R90_512x8m81_1
timestamp 1763476864
transform 0 -1 333 1 0 11621
box 0 0 65 89
<< labels >>
rlabel metal1 s 229 10312 229 10312 4 pcb
port 8 nsew
rlabel metal3 s 303 6306 303 6306 4 vss
port 1 nsew
rlabel metal3 s 318 11384 318 11384 4 vdd
port 2 nsew
rlabel metal2 s 125 11421 125 11421 4 bb
port 4 nsew
rlabel metal2 s 441 11421 441 11421 4 b
port 3 nsew
rlabel metal2 s 54 3775 54 3775 4 db
port 5 nsew
rlabel metal2 s 44 3775 44 3775 6 db
port 5 nsew
rlabel metal1 s 318 4597 318 4597 4 vdd
port 2 nsew
rlabel metal2 s 261 4463 261 4463 4 ypass
port 6 nsew
<< properties >>
string path 0.000 27.385 0.000 -0.005 
<< end >>
