magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nwell >>
rect -78 150 771 835
rect -78 -189 637 150
<< pmos >>
rect 96 236 597 749
<< pdiff >>
rect 8 736 96 749
rect 8 249 21 736
rect 67 249 96 736
rect 8 236 96 249
rect 597 735 685 749
rect 597 249 626 735
rect 672 249 685 735
rect 597 236 685 249
<< pdiffc >>
rect 21 249 67 736
rect 626 249 672 735
<< psubdiff >>
rect 8 928 670 1001
<< nsubdiff >>
rect 38 36 520 138
<< polysilicon >>
rect 96 749 597 843
rect 96 191 597 236
<< metal1 >>
rect 0 966 678 1001
rect 0 810 2 966
rect 58 810 678 966
rect 0 795 678 810
rect 9 736 100 739
rect 9 249 21 736
rect 67 249 100 736
rect 9 240 100 249
rect 592 735 683 739
rect 592 249 626 735
rect 672 249 683 735
rect 592 240 683 249
rect 38 36 520 138
<< via1 >>
rect 2 810 58 966
<< metal2 >>
rect 0 966 60 983
rect 0 810 2 966
rect 58 810 60 966
rect 0 795 60 810
rect 22 240 670 651
<< via2 >>
rect 2 810 58 966
<< metal3 >>
rect -2 966 92 1517
rect -2 810 2 966
rect 58 810 106 966
rect -2 0 92 810
rect 307 0 401 1028
rect 600 0 694 1028
use M1_NACTIVE_01_R270_3v256x8m81  M1_NACTIVE_01_R270_3v256x8m81_0
timestamp 1763766357
transform 1 0 282 0 1 102
box -284 -54 284 53
use M1_PACTIVE_R270_3v256x8m81  M1_PACTIVE_R270_3v256x8m81_0
timestamp 1763766357
transform 1 0 342 0 1 964
box -284 -36 284 37
use M1_POLY2_01_R270_3v256x8m81  M1_POLY2_01_R270_3v256x8m81_0
timestamp 1763766357
transform 1 0 350 0 1 821
box -240 -46 240 46
use M2_M1$04_R270_3v256x8m81  M2_M1$04_R270_3v256x8m81_0
timestamp 1763766357
transform 1 0 41 0 1 465
box -46 -266 46 266
<< end >>
