magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< nwell >>
rect -202 -86 362 437
<< pmos >>
rect -28 0 28 351
rect 132 0 188 351
<< pdiff >>
rect -116 338 -28 351
rect -116 13 -103 338
rect -57 13 -28 338
rect -116 0 -28 13
rect 28 338 132 351
rect 28 13 57 338
rect 103 13 132 338
rect 28 0 132 13
rect 188 338 276 351
rect 188 13 217 338
rect 263 13 276 338
rect 188 0 276 13
<< pdiffc >>
rect -103 13 -57 338
rect 57 13 103 338
rect 217 13 263 338
<< polysilicon >>
rect -28 351 28 395
rect 132 351 188 395
rect -28 -44 28 0
rect 132 -44 188 0
<< metal1 >>
rect -103 338 -57 351
rect -103 0 -57 13
rect 57 338 103 351
rect 57 0 103 13
rect 217 338 263 351
rect 217 0 263 13
<< labels >>
flabel pdiffc 80 175 80 175 0 FreeSans 186 0 0 0 D
flabel pdiffc -68 175 -68 175 0 FreeSans 186 0 0 0 S
flabel pdiffc 228 175 228 175 0 FreeSans 186 0 0 0 S
<< end >>
