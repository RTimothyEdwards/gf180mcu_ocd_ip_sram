magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -119 476 119 511
rect -119 -781 -93 476
rect 93 -781 119 476
rect -119 -808 119 -781
<< via2 >>
rect -93 -781 93 476
<< metal3 >>
rect -119 476 119 511
rect -119 -781 -93 476
rect 93 -781 119 476
rect -119 -808 119 -781
<< end >>
