magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< error_p >>
rect -45 -297 -44 -285
rect 44 -297 45 -285
<< metal1 >>
rect -40 959 39 961
rect -44 940 44 959
rect -44 -297 -26 940
rect -45 -310 -26 -297
rect 26 -297 44 940
rect 26 -310 45 -297
rect -45 -331 45 -310
<< via1 >>
rect -26 -310 26 940
<< metal2 >>
rect -44 940 44 959
rect -44 -310 -26 940
rect 26 -310 44 940
rect -44 -331 44 -310
<< end >>
