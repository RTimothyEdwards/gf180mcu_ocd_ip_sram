magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal1 >>
rect -113 235 113 243
rect -113 -235 -105 235
rect 105 -235 113 235
rect -113 -243 113 -235
<< via1 >>
rect -105 -235 105 235
<< metal2 >>
rect -113 235 113 243
rect -113 -235 -105 235
rect 105 -235 113 235
rect -113 -243 113 -235
<< end >>
