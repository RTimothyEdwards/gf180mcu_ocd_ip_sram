magic
tech gf180mcuD
magscale 1 10
timestamp 1765833632
<< nwell >>
rect 120 5529 1129 5843
rect 295 3977 299 5529
rect 854 3977 1000 5529
<< nmos >>
rect 483 2025 539 3169
rect 612 2025 668 3169
<< ndiff >>
rect 373 3145 483 3169
rect 373 2137 396 3145
rect 442 2137 483 3145
rect 373 2025 483 2137
rect 539 2025 612 3169
rect 668 3144 779 3169
rect 668 2137 710 3144
rect 756 2137 779 3144
rect 668 2025 779 2137
<< ndiffc >>
rect 396 2137 442 3145
rect 710 2137 756 3144
<< psubdiff >>
rect 889 3134 982 3169
rect 889 1973 911 3134
rect 959 1973 982 3134
rect 889 1938 982 1973
rect 288 1913 1009 1938
rect 288 1867 338 1913
rect 847 1867 1009 1913
rect 288 1842 1009 1867
<< nsubdiff >>
rect 206 5694 1043 5727
rect 206 5648 320 5694
rect 436 5648 720 5694
rect 867 5648 1043 5694
rect 206 5615 1043 5648
<< psubdiffcont >>
rect 911 1973 959 3134
rect 338 1867 847 1913
<< nsubdiffcont >>
rect 320 5648 436 5694
rect 720 5648 867 5694
<< polysilicon >>
rect 347 7117 403 7265
rect 507 7117 563 7265
rect 667 7117 723 7265
rect 827 7117 883 7265
rect 347 7044 883 7117
rect 347 7027 403 7044
rect 507 7027 563 7044
rect 667 7027 723 7044
rect 827 7027 883 7044
rect 347 5883 403 5891
rect 507 5883 563 5891
rect 667 5883 723 5891
rect 827 5883 883 5891
rect 345 5788 899 5883
rect 472 3984 528 4037
rect 472 3898 539 3984
rect 483 3169 539 3898
rect 632 3743 688 4037
rect 612 3675 688 3743
rect 612 3169 668 3675
rect 483 1974 539 2025
rect 612 1974 668 2025
<< metal1 >>
rect 268 7980 932 7982
rect 268 7922 976 7980
rect 268 7646 349 7922
rect 581 7646 662 7922
rect 895 7646 976 7922
rect 416 7125 498 7366
rect 738 7125 819 7216
rect 416 7041 819 7125
rect 416 6936 498 7041
rect 738 6936 819 7041
rect 346 5794 898 5877
rect 535 5793 617 5794
rect 170 5694 459 5712
rect 170 5648 320 5694
rect 436 5648 459 5694
rect 170 5629 459 5648
rect 378 5628 459 5629
rect 378 5556 460 5628
rect 535 4058 616 5793
rect 692 5694 1043 5712
rect 692 5648 720 5694
rect 867 5648 1043 5694
rect 692 5629 1043 5648
rect 692 4069 976 5629
rect 255 3901 1068 3965
rect 255 3759 1068 3824
rect 255 3619 1068 3683
rect 255 3263 1068 3542
rect 378 3145 459 3162
rect 378 2137 396 3145
rect 442 2137 459 3145
rect 378 2031 459 2137
rect 692 3144 976 3162
rect 692 2137 710 3144
rect 756 3134 976 3144
rect 756 2137 911 3134
rect 692 1973 911 2137
rect 959 1973 976 3134
rect 692 1942 976 1973
rect 692 1935 981 1942
rect 288 1913 1009 1935
rect 288 1867 338 1913
rect 847 1867 1009 1913
rect 288 1845 1009 1867
<< metal2 >>
rect 734 7187 889 7809
rect 692 4902 981 5678
rect 374 4069 620 4314
rect 374 2920 464 4069
rect 692 1783 981 3162
<< metal3 >>
rect 107 7657 1038 7758
rect 107 7179 1039 7657
rect 107 6575 1038 7043
rect 107 5938 1036 6500
rect 107 4362 1036 5857
rect 598 2766 1038 3243
rect 598 2319 1039 2682
rect 598 1785 1041 2247
use M1_NACTIVE4310591302024_3v256x8m81  M1_NACTIVE4310591302024_3v256x8m81_0
timestamp 1765833244
transform 1 0 936 0 1 4275
box -38 -128 36 128
use M1_POLY24310591302059_3v256x8m81  M1_POLY24310591302059_3v256x8m81_0
timestamp 1763766357
transform 1 0 605 0 1 5835
box -161 -36 161 36
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_0
timestamp 1765833244
transform -1 0 576 0 1 4192
box -43 -122 43 122
use M2_M1$$43376684_3v256x8m81  M2_M1$$43376684_3v256x8m81_0
timestamp 1763766357
transform -1 0 419 0 1 2583
box -44 21 44 579
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_0
timestamp 1763766357
transform 1 0 779 0 1 7462
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_1
timestamp 1763766357
transform 1 0 616 0 1 7462
box -44 -275 44 275
use M2_M1$$43379756_3v256x8m81  M2_M1$$43379756_3v256x8m81_2
timestamp 1763766357
transform -1 0 295 0 1 7462
box -44 -275 44 275
use M2_M1$$43380780_3v256x8m81  M2_M1$$43380780_3v256x8m81_0
timestamp 1763766357
transform -1 0 295 0 1 6775
box -44 -198 44 198
use M2_M1$$43380780_3v256x8m81  M2_M1$$43380780_3v256x8m81_1
timestamp 1763766357
transform 1 0 622 0 1 6775
box -44 -198 44 198
use M2_M1$$43380780_3v256x8m81  M2_M1$$43380780_3v256x8m81_2
timestamp 1763766357
transform 1 0 935 0 1 6775
box -44 -198 44 198
use M2_M1$$47500332_3v256x8m81  M2_M1$$47500332_3v256x8m81_0
timestamp 1763766357
transform 1 0 737 0 1 4835
box -44 -432 44 732
use M2_M1$$47500332_3v256x8m81  M2_M1$$47500332_3v256x8m81_1
timestamp 1763766357
transform 1 0 421 0 1 4835
box -44 -432 44 732
use M2_M1$$47500332_3v256x8m81  M2_M1$$47500332_3v256x8m81_2
timestamp 1763766357
transform 1 0 935 0 1 4835
box -44 -432 44 732
use M2_M1$$47640620_3v256x8m81  M2_M1$$47640620_3v256x8m81_0
timestamp 1763766357
transform 1 0 935 0 1 2182
box -45 -84 45 884
use M2_M1$$47640620_3v256x8m81  M2_M1$$47640620_3v256x8m81_1
timestamp 1763766357
transform 1 0 737 0 1 2182
box -45 -84 45 884
use M3_M2$$47108140_3v256x8m81  M3_M2$$47108140_3v256x8m81_0
timestamp 1763766357
transform 1 0 935 0 1 2967
box -45 -198 45 198
use M3_M2$$47108140_3v256x8m81  M3_M2$$47108140_3v256x8m81_1
timestamp 1763766357
transform 1 0 737 0 1 2967
box -45 -198 45 198
use M3_M2$$47108140_3v256x8m81  M3_M2$$47108140_3v256x8m81_2
timestamp 1763766357
transform -1 0 295 0 1 6785
box -45 -198 45 198
use M3_M2$$47108140_3v256x8m81  M3_M2$$47108140_3v256x8m81_3
timestamp 1763766357
transform 1 0 622 0 1 6785
box -45 -198 45 198
use M3_M2$$47108140_3v256x8m81  M3_M2$$47108140_3v256x8m81_4
timestamp 1763766357
transform 1 0 935 0 1 6785
box -45 -198 45 198
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_0
timestamp 1763766357
transform 1 0 935 0 1 1970
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_1
timestamp 1763766357
transform 1 0 737 0 1 1970
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_2
timestamp 1763766357
transform 1 0 616 0 1 7462
box -84 -185 84 275
use M3_M2$$47333420_3v256x8m81  M3_M2$$47333420_3v256x8m81_3
timestamp 1763766357
transform -1 0 295 0 1 7462
box -84 -185 84 275
use M3_M2$$47644716_3v256x8m81  M3_M2$$47644716_3v256x8m81_0
timestamp 1763766357
transform 1 0 737 0 1 4835
box -45 -432 45 732
use M3_M2$$47644716_3v256x8m81  M3_M2$$47644716_3v256x8m81_1
timestamp 1763766357
transform 1 0 421 0 1 4835
box -45 -432 45 732
use M3_M2$$47644716_3v256x8m81  M3_M2$$47644716_3v256x8m81_2
timestamp 1763766357
transform 1 0 935 0 1 4835
box -45 -432 45 732
use nmos_1p2$$47641644_3v256x8m81  nmos_1p2$$47641644_3v256x8m81_0
timestamp 1763766357
transform -1 0 869 0 -1 7726
box -102 -44 130 467
use nmos_1p2$$47641644_3v256x8m81  nmos_1p2$$47641644_3v256x8m81_1
timestamp 1763766357
transform -1 0 549 0 -1 7726
box -102 -44 130 467
use nmos_1p2$$47641644_3v256x8m81  nmos_1p2$$47641644_3v256x8m81_2
timestamp 1763766357
transform -1 0 389 0 -1 7726
box -102 -44 130 467
use nmos_1p2$$47641644_3v256x8m81  nmos_1p2$$47641644_3v256x8m81_3
timestamp 1763766357
transform -1 0 709 0 -1 7726
box -102 -44 130 467
use pmos_1p2$$47513644_3v256x8m81  pmos_1p2$$47513644_3v256x8m81_0
timestamp 1763766357
transform -1 0 709 0 -1 6985
box -188 -86 216 1144
use pmos_1p2$$47513644_3v256x8m81  pmos_1p2$$47513644_3v256x8m81_1
timestamp 1763766357
transform -1 0 549 0 -1 6985
box -188 -86 216 1144
use pmos_1p2$$47513644_3v256x8m81  pmos_1p2$$47513644_3v256x8m81_2
timestamp 1763766357
transform -1 0 389 0 -1 6985
box -188 -86 216 1144
use pmos_1p2$$47513644_3v256x8m81  pmos_1p2$$47513644_3v256x8m81_3
timestamp 1763766357
transform -1 0 869 0 -1 6985
box -188 -86 216 1144
use pmos_1p2$$47642668_3v256x8m81  pmos_1p2$$47642668_3v256x8m81_0
timestamp 1763766357
transform -1 0 674 0 1 4063
box -194 -86 220 1504
use pmos_1p2$$47643692_3v256x8m81  pmos_1p2$$47643692_3v256x8m81_0
timestamp 1763766357
transform -1 0 514 0 1 4063
box -188 -86 216 1504
<< end >>
