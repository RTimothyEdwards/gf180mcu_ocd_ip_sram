magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal1 >>
rect -783 26 783 46
rect -783 -26 -764 26
rect 764 -26 783 26
rect -783 -46 783 -26
<< via1 >>
rect -764 -26 764 26
<< metal2 >>
rect -782 26 783 46
rect -782 -26 -764 26
rect 764 -26 783 26
rect -782 -46 783 -26
<< end >>
