magic
tech gf180mcuD
magscale 1 10
timestamp 1766784746
<< nwell >>
rect 8121 20390 8391 20405
rect 939 17073 15865 20390
rect 15938 20389 16273 20408
rect 851 13113 15617 13972
rect 15636 13226 16048 13972
rect 15636 13113 16208 13226
rect 15899 13112 16208 13113
rect 15905 13110 16208 13112
rect 15978 10713 16689 11141
rect 16016 6294 16103 6426
rect 4187 6217 4464 6269
rect 12056 6220 12118 6237
<< metal1 >>
rect 359 20805 523 21208
rect 4267 20816 4431 21206
rect 8175 20813 8339 21209
rect 12083 20815 12247 21203
rect 15989 20873 16153 21205
rect 15989 20754 17384 20873
rect 15584 18915 16039 18973
rect 16364 13783 16606 14445
rect 664 -470 898 -410
<< metal2 >>
rect 253 20629 323 21827
rect 555 19283 625 21827
rect 8063 20661 8133 21827
rect 8365 19268 8435 21827
rect 15873 19268 15943 21827
rect 16195 20706 16265 21827
rect 16155 20629 16265 20706
rect 16155 19268 16225 20629
rect 675 1791 740 1991
rect 1293 1786 1359 1986
rect 7347 1909 7413 2109
rect 7959 1909 8024 2109
rect 8491 1792 8556 1992
rect 9109 1787 9175 1987
rect 15163 1910 15229 2110
rect 15775 1910 15840 2110
<< metal3 >>
rect 0 41725 16576 41865
rect 0 21475 16576 21727
rect -367 21117 16576 21274
rect 0 20661 16860 20997
rect 560 19107 16860 20373
rect 722 15512 15882 15662
rect 722 15511 921 15512
rect 722 15266 15882 15418
rect 722 15022 15882 15172
rect 722 14776 15882 14927
rect 724 14553 15882 14704
rect 724 14312 15882 14463
rect 724 14062 15882 14212
rect 724 13818 15882 13969
rect 919 13362 15920 13672
rect 919 12774 15920 13094
rect 927 11344 16276 11944
rect 919 10037 16276 11344
rect 919 7981 16276 9834
rect 883 7355 16597 7856
rect 883 6419 17141 6986
rect 919 5118 16779 6042
rect 815 4957 15796 5018
rect 815 4774 16513 4841
rect 919 3704 16916 4657
rect 919 3121 16993 3483
rect 919 3044 16276 3064
rect 529 2718 16276 3044
rect 919 2353 16862 2656
rect 919 1941 17155 2260
rect 893 1234 17221 1553
rect 893 786 16276 1033
rect 893 477 16276 538
rect 893 144 16274 390
rect 893 -196 16276 -45
rect 893 -364 16274 -196
use dcap_103_novia_3v256x8m81  dcap_103_novia_3v256x8m81_0
array 0 35 452 0 0 552
timestamp 1765833244
transform 1 0 -39 0 1 20404
box -205 -132 492 420
use M2_M1$$43374636_3v256x8m81  M2_M1$$43374636_3v256x8m81_0
timestamp 1765833244
transform 1 0 16400 0 1 4856
box -119 -123 119 123
use M2_M1431059130200_3v256x8m81  M2_M1431059130200_3v256x8m81_0
timestamp 1765833244
transform -1 0 16192 0 -1 20811
box -63 -34 63 34
use M2_M1431059130200_3v256x8m81  M2_M1431059130200_3v256x8m81_1
timestamp 1765833244
transform -1 0 8099 0 -1 20784
box -63 -34 63 34
use M2_M1431059130200_3v256x8m81  M2_M1431059130200_3v256x8m81_2
timestamp 1765833244
transform -1 0 294 0 -1 20785
box -63 -34 63 34
use M3_M2$$201416748_3v256x8m81  M3_M2$$201416748_3v256x8m81_0
timestamp 1765833244
transform 1 0 16400 0 1 4859
box -119 -123 119 123
use M3_M24310591302022_3v256x8m81  M3_M24310591302022_3v256x8m81_0
timestamp 1765833244
transform 1 0 8400 0 1 19821
box -35 -534 35 534
use M3_M24310591302022_3v256x8m81  M3_M24310591302022_3v256x8m81_1
timestamp 1765833244
transform 1 0 15908 0 1 19821
box -35 -534 35 534
use M3_M24310591302022_3v256x8m81  M3_M24310591302022_3v256x8m81_2
timestamp 1765833244
transform 1 0 590 0 1 19821
box -35 -534 35 534
use M3_M24310591302023_3v256x8m81  M3_M24310591302023_3v256x8m81_0
timestamp 1765833244
transform 1 0 286 0 1 20832
box -35 -165 35 165
use M3_M24310591302023_3v256x8m81  M3_M24310591302023_3v256x8m81_1
timestamp 1765833244
transform 1 0 8098 0 1 20832
box -35 -165 35 165
use M3_M24310591302023_3v256x8m81  M3_M24310591302023_3v256x8m81_2
timestamp 1765833244
transform 1 0 16230 0 1 20832
box -35 -165 35 165
use rarray4_256_3v256x8m81  rarray4_256_3v256x8m81_0
timestamp 1765833452
transform 1 0 321 0 1 21628
box -1397 103 16315 19939
use rdummy_3v256x4_3v256x8m81  rdummy_3v256x4_3v256x8m81_0
timestamp 1765981949
transform 1 0 214 0 1 21064
box -631 -16314 16729 20854
use saout_m2_3v256x8m81  saout_m2_3v256x8m81_2
timestamp 1766784746
transform 1 0 8164 0 1 0
box -188 -475 5343 21797
use saout_m2_3v256x8m81  saout_m2_3v256x8m81_3
timestamp 1766784746
transform 1 0 348 0 1 -1
box -188 -475 5343 21797
use saout_R_m2_3v256x8m81  saout_R_m2_3v256x8m81_1
timestamp 1766784746
transform -1 0 16164 0 1 5
box -188 -482 5343 21793
use saout_R_m2_3v256x8m81  saout_R_m2_3v256x8m81_3
timestamp 1766784746
transform -1 0 8348 0 1 4
box -188 -482 5343 21793
<< labels >>
rlabel metal3 s 1125 40367 1125 40367 4 WL[29]
port 21 nsew
rlabel metal3 s 1125 37847 1125 37847 4 WL[25]
port 22 nsew
rlabel metal3 s 1125 37217 1125 37217 4 WL[24]
port 23 nsew
rlabel metal3 s 1125 36587 1125 36587 4 WL[23]
port 24 nsew
rlabel metal3 s 1125 35957 1125 35957 4 WL[22]
port 25 nsew
rlabel metal3 s 1125 34697 1125 34697 4 WL[20]
port 26 nsew
rlabel metal3 s 1125 39107 1125 39107 4 WL[27]
port 27 nsew
rlabel metal3 s 1125 40997 1125 40997 4 WL[30]
port 28 nsew
rlabel metal3 s 1125 33437 1125 33437 4 WL[18]
port 29 nsew
rlabel metal3 s 1125 31547 1125 31547 4 WL[15]
port 31 nsew
rlabel metal3 s 1125 41627 1125 41627 4 WL[31]
port 37 nsew
rlabel metal3 s 1125 30917 1125 30917 4 WL[14]
port 38 nsew
rlabel metal3 s 1125 32177 1125 32177 4 WL[16]
port 39 nsew
rlabel metal3 s 1125 32807 1125 32807 4 WL[17]
port 40 nsew
rlabel metal3 s 1125 38477 1125 38477 4 WL[26]
port 41 nsew
rlabel metal3 s 1125 34067 1125 34067 4 WL[19]
port 42 nsew
rlabel metal3 s 1125 39737 1125 39737 4 WL[28]
port 46 nsew
rlabel metal3 s 1125 35327 1125 35327 4 WL[21]
port 48 nsew
rlabel metal3 s 1125 22097 1125 22097 4 WL[0]
port 53 nsew
rlabel metal3 s 1125 23357 1125 23357 4 WL[2]
port 54 nsew
rlabel metal3 s 1125 29657 1125 29657 4 WL[12]
port 55 nsew
rlabel metal3 s 1125 23987 1125 23987 4 WL[3]
port 56 nsew
rlabel metal3 s 1125 24617 1125 24617 4 WL[4]
port 57 nsew
rlabel metal3 s 1125 26507 1125 26507 4 WL[7]
port 59 nsew
rlabel metal3 s 1125 27137 1125 27137 4 WL[8]
port 60 nsew
rlabel metal3 s 1125 27767 1125 27767 4 WL[9]
port 61 nsew
rlabel metal3 s 1125 22727 1125 22727 4 WL[1]
port 62 nsew
rlabel metal3 s 1124 25247 1124 25247 4 WL[5]
port 65 nsew
rlabel metal3 s 1125 28397 1125 28397 4 WL[10]
port 67 nsew
rlabel metal3 s 1125 30287 1125 30287 4 WL[13]
port 68 nsew
rlabel metal3 s 1124 25877 1124 25877 4 WL[6]
port 75 nsew
rlabel metal3 s 1125 29027 1125 29027 4 WL[11]
port 79 nsew
rlabel metal3 s 168 21213 168 21213 4 VSS
port 18 nsew
rlabel metal3 s 942 4999 942 4999 4 GWE
port 78 nsew
rlabel metal3 s 942 4819 942 4819 4 tblhl
port 76 nsew
flabel metal1 s 15725 -438 15725 -438 0 FreeSans 420 0 0 0 WEN[4]
port 92 nsew
flabel metal1 s 8650 -438 8650 -438 0 FreeSans 420 0 0 0 WEN[5]
port 95 nsew
flabel metal1 s 7950 -438 7950 -438 0 FreeSans 420 0 0 0 WEN[6]
port 96 nsew
flabel metal1 s 693 -446 693 -446 0 FreeSans 420 0 0 0 WEN[7]
port 93 nsew
rlabel metal2 s 1319 1882 1319 1882 4 q[4]
port 87 nsew
rlabel metal2 s 700 1830 700 1830 4 din[4]
port 97 se
rlabel metal2 s 7372 1926 7372 1926 4 q[5]
port 82 nsew
rlabel metal2 s 7990 1922 7990 1922 4 din[5]
port 85 nsew
rlabel metal2 s 8527 1822 8527 1822 4 din[6]
port 86 nsew
rlabel metal2 s 9141 1882 9141 1882 4 q[6]
port 83 nsew
rlabel metal2 s 15183 1922 15183 1922 4 q[7]
port 84 nsew
rlabel metal2 s 15814 1922 15814 1922 4 din[7]
port 81 nsew
rlabel metal3 780 19700 780 19700 4 VDD
port 98 se
rlabel metal3 4320 -230 4320 -230 0 VDD
rlabel metal3 4210 1380 4210 1380 0 VDD
rlabel metal3 4180 2090 4180 2090 0 VDD
rlabel metal3 4260 4200 4260 4200 0 VDD
rlabel metal3 4350 6710 4350 6710 0 VDD
rlabel metal3 4290 10760 4290 10760 0 VDD
rlabel metal3 4230 13510 4230 13510 0 VDD
rlabel metal1 s 3184 11809 3184 11809 4 pcb[7]
port 89 nsew
rlabel metal1 s 5489 11789 5489 11789 4 pcb[6]
port 88 nsew
rlabel metal1 s 11001 11799 11001 11799 4 pcb[5]
port 94 nsew
rlabel metal1 s 13306 11799 13306 11799 4 pcb[4]
port 90 nsew
<< end >>
