magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -70 106 70 113
rect -70 -106 -63 106
rect 63 -106 70 106
rect -70 -113 70 -106
<< via2 >>
rect -63 -106 63 106
<< metal3 >>
rect -70 106 70 113
rect -70 -106 -63 106
rect 63 -106 70 106
rect -70 -113 70 -106
<< end >>
