magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< polysilicon >>
rect -96 211 -41 245
rect 63 211 119 245
rect 223 211 279 245
rect 383 211 439 245
rect -96 -34 -41 0
rect 63 -34 119 0
rect 223 -34 279 0
rect 383 -34 439 0
use nmos_5p04310591302012_3v512x8m81  nmos_5p04310591302012_3v512x8m81_0
timestamp 1764525316
transform 1 0 -14 0 1 0
box -171 -44 541 255
<< end >>
