magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< nwell >>
rect -133 -66 265 383
<< polysilicon >>
rect -42 317 13 351
rect 118 317 173 351
rect -42 -34 13 0
rect 118 -34 174 0
use pmos_5p04310591302031_512x8m81  pmos_5p04310591302031_512x8m81_0
timestamp 1763765945
transform 1 0 -14 0 1 0
box -202 -86 362 404
<< end >>
