magic
tech gf180mcuD
magscale 1 10
timestamp 1765213032
<< nwell >>
rect -133 1589 3403 2104
rect 941 485 1137 487
rect -133 0 3403 485
<< pdiff >>
rect 1205 1687 1287 1822
rect 1458 1687 1498 1822
<< polysilicon >>
rect 253 1936 309 2049
rect 737 2039 1370 2062
rect 737 2006 1371 2039
rect 737 1931 793 2006
rect 1315 1817 1371 2006
rect 253 1409 309 1651
rect 413 1409 469 1651
rect 737 1636 793 1651
rect 716 1564 793 1636
rect 869 1595 1138 1644
rect 869 1587 1459 1595
rect 737 1432 793 1564
rect 1076 1539 1459 1587
rect 1403 1484 1459 1539
rect 1563 1563 1625 1662
rect 1563 1489 1619 1563
rect 1873 1478 1929 1659
rect 2033 1478 2089 1659
rect 2346 1597 2402 1732
rect 2501 1597 2557 1732
rect 2819 1597 2875 1648
rect 2979 1597 3035 1648
rect 2346 1560 3195 1597
rect 2350 1556 3195 1560
rect 2501 1456 2557 1556
rect 3139 1417 3195 1556
rect 413 1155 469 1213
rect 737 1131 793 1271
rect 1873 1189 1929 1333
rect 1701 1133 1929 1189
rect 2033 1132 2089 1323
rect 737 1075 1135 1131
rect 2819 1120 2875 1139
rect 2979 1120 3035 1139
rect 2561 1101 3035 1120
rect 2561 1079 3033 1101
rect 419 882 475 953
rect 1258 823 1314 903
rect 259 440 315 717
rect 419 440 475 717
rect 737 559 793 670
rect 712 487 793 559
rect 737 437 793 487
rect 1260 532 1316 619
rect 1794 551 1850 674
rect 1954 551 2010 674
rect 2115 551 2171 674
rect 1260 491 1477 532
rect 1794 500 2171 551
rect 1260 437 1316 491
rect 1420 440 1476 491
rect 1794 441 1850 500
rect 1954 441 2010 500
rect 2115 441 2171 500
rect 259 23 315 153
<< metal1 >>
rect 212 2207 2971 2300
rect 212 2058 325 2207
rect 165 1694 256 2005
rect 483 1631 564 2005
rect 635 1694 725 2005
rect 326 1572 698 1631
rect 326 1246 407 1572
rect 792 1304 882 2005
rect 479 1096 569 1272
rect 991 1110 1080 2005
rect 1148 1822 1237 2005
rect 1487 1822 1534 1895
rect 1148 1687 1294 1822
rect 1419 1687 1534 1822
rect 1626 1694 1717 2005
rect 1148 1492 1237 1687
rect 1148 1358 1399 1492
rect 1487 1435 1534 1687
rect 1784 1632 1873 2005
rect 1940 1694 2031 2005
rect 1723 1566 1873 1632
rect 1500 1358 1532 1435
rect 1148 1192 1237 1358
rect 1784 1192 1873 1566
rect 2097 1619 2187 2005
rect 2097 1571 2352 1619
rect 2097 1358 2187 1571
rect 1148 1144 1717 1192
rect 1784 1144 2147 1192
rect 821 1060 1080 1110
rect 2411 1091 2501 2006
rect 2725 1631 2814 2005
rect 2881 1694 2971 2207
rect 3038 1631 3128 2005
rect 2725 1547 3128 1631
rect 351 760 383 767
rect 343 554 391 760
rect 343 506 631 554
rect 165 92 256 401
rect 502 373 550 506
rect 634 84 725 401
rect 821 324 871 1060
rect 2725 1034 2814 1547
rect 2881 1173 2972 1485
rect 3038 1034 3128 1547
rect 3194 1173 3285 1491
rect 1268 980 3128 1034
rect 1275 900 1307 980
rect 1344 555 1397 701
rect 1344 539 1777 555
rect 1879 549 1927 774
rect 2198 549 2245 790
rect 1344 507 1780 539
rect 1344 498 1777 507
rect 1166 84 1257 401
rect 1344 376 1397 498
rect 1879 465 2531 549
rect 1480 84 1571 401
rect 1698 84 1789 401
rect 1879 376 1927 465
rect 2012 84 2103 401
rect 2198 376 2245 465
rect 91 -16 325 36
<< metal2 >>
rect 991 1179 1080 2005
rect 2881 1179 2972 2004
<< metal3 >>
rect -45 1687 3403 2006
rect -45 1240 3403 1486
rect -45 1092 3403 1153
rect -45 930 3403 991
rect -45 597 3403 842
rect -45 89 3403 408
use M1_NACTIVE4310591302037_3v1024x8m81  M1_NACTIVE4310591302037_3v1024x8m81_0
timestamp 1764692000
transform 1 0 2594 0 1 273
box -135 -158 135 158
use M1_NACTIVE_01_3v1024x8m81  M1_NACTIVE_01_3v1024x8m81_0
timestamp 1764692000
transform 1 0 2380 0 1 256
box -139 -198 139 199
use M1_NACTIVE_01_3v1024x8m81  M1_NACTIVE_01_3v1024x8m81_1
timestamp 1764692000
transform 1 0 1026 0 1 256
box -139 -198 139 199
use M1_NACTIVE_01_3v1024x8m81  M1_NACTIVE_01_3v1024x8m81_2
timestamp 1764692000
transform 1 0 0 0 1 256
box -139 -198 139 199
use M1_NACTIVE_01_3v1024x8m81  M1_NACTIVE_01_3v1024x8m81_3
timestamp 1764692000
transform 1 0 0 0 1 1854
box -139 -198 139 199
use M1_NACTIVE_01_3v1024x8m81  M1_NACTIVE_01_3v1024x8m81_4
timestamp 1764692000
transform 1 0 3294 0 1 1854
box -139 -198 139 199
use M1_PACTIVE4310591302027_3v1024x8m81  M1_PACTIVE4310591302027_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2380 0 1 716
box -53 -62 53 62
use M1_PACTIVE4310591302027_3v1024x8m81  M1_PACTIVE4310591302027_3v1024x8m81_1
timestamp 1764525316
transform 1 0 2 0 1 716
box -53 -62 53 62
use M1_PACTIVE4310591302027_3v1024x8m81  M1_PACTIVE4310591302027_3v1024x8m81_2
timestamp 1764525316
transform 1 0 1024 0 1 716
box -53 -62 53 62
use M1_PACTIVE4310591302027_3v1024x8m81  M1_PACTIVE4310591302027_3v1024x8m81_3
timestamp 1764525316
transform 1 0 1530 0 1 716
box -53 -62 53 62
use M1_PACTIVE4310591302027_3v1024x8m81  M1_PACTIVE4310591302027_3v1024x8m81_4
timestamp 1764525316
transform 1 0 2 0 1 1365
box -53 -62 53 62
use M1_PACTIVE4310591302027_3v1024x8m81  M1_PACTIVE4310591302027_3v1024x8m81_5
timestamp 1764525316
transform 1 0 3418 0 1 1365
box -53 -62 53 62
use M1_POLY24310591302019_3v1024x8m81  M1_POLY24310591302019_3v1024x8m81_0
timestamp 1764525316
transform 0 -1 644 -1 0 1600
box -36 -80 36 78
use M1_POLY24310591302019_3v1024x8m81  M1_POLY24310591302019_3v1024x8m81_1
timestamp 1764525316
transform 1 0 906 0 1 1542
box -36 -80 36 78
use M1_POLY24310591302019_3v1024x8m81  M1_POLY24310591302019_3v1024x8m81_2
timestamp 1764525316
transform 0 -1 2301 1 0 1595
box -36 -80 36 78
use M1_POLY24310591302019_3v1024x8m81  M1_POLY24310591302019_3v1024x8m81_3
timestamp 1764525316
transform 0 -1 2135 1 0 1168
box -36 -80 36 78
use M1_POLY24310591302019_3v1024x8m81  M1_POLY24310591302019_3v1024x8m81_4
timestamp 1764525316
transform 0 -1 2500 1 0 1115
box -36 -80 36 78
use M1_POLY24310591302019_3v1024x8m81  M1_POLY24310591302019_3v1024x8m81_5
timestamp 1764525316
transform 0 -1 1684 1 0 1596
box -36 -80 36 78
use M1_POLY24310591302019_3v1024x8m81  M1_POLY24310591302019_3v1024x8m81_6
timestamp 1764525316
transform 0 -1 1652 1 0 1168
box -36 -80 36 78
use M1_POLY24310591302033_3v1024x8m81  M1_POLY24310591302033_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1747 0 1 523
box -62 -36 62 36
use M1_POLY24310591302033_3v1024x8m81  M1_POLY24310591302033_3v1024x8m81_1
timestamp 1764525316
transform 0 -1 1291 1 0 955
box -62 -36 62 36
use M1_POLY24310591302033_3v1024x8m81  M1_POLY24310591302033_3v1024x8m81_2
timestamp 1764525316
transform 1 0 268 0 1 12
box -62 -36 62 36
use M1_POLY24310591302033_3v1024x8m81  M1_POLY24310591302033_3v1024x8m81_3
timestamp 1764525316
transform 1 0 466 0 1 961
box -62 -36 62 36
use M1_POLY24310591302033_3v1024x8m81  M1_POLY24310591302033_3v1024x8m81_4
timestamp 1764525316
transform 1 0 655 0 1 523
box -62 -36 62 36
use M1_POLY24310591302033_3v1024x8m81  M1_POLY24310591302033_3v1024x8m81_5
timestamp 1764525316
transform 1 0 466 0 1 1123
box -62 -36 62 36
use M1_POLY24310591302033_3v1024x8m81  M1_POLY24310591302033_3v1024x8m81_6
timestamp 1764525316
transform 1 0 268 0 1 2082
box -62 -36 62 36
use M2_M1$$202395692_3v1024x8m81  M2_M1$$202395692_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2058 0 1 256
box -44 -111 44 112
use M2_M1$$202395692_3v1024x8m81  M2_M1$$202395692_3v1024x8m81_1
timestamp 1764525316
transform 1 0 1744 0 1 730
box -44 -111 44 112
use M2_M1$$202395692_3v1024x8m81  M2_M1$$202395692_3v1024x8m81_2
timestamp 1764525316
transform 1 0 1744 0 1 256
box -44 -111 44 112
use M2_M1$$202395692_3v1024x8m81  M2_M1$$202395692_3v1024x8m81_3
timestamp 1764525316
transform 1 0 2058 0 1 730
box -44 -111 44 112
use M2_M1$$202395692_3v1024x8m81  M2_M1$$202395692_3v1024x8m81_4
timestamp 1764525316
transform 1 0 524 0 1 730
box -44 -111 44 112
use M2_M1$$202395692_3v1024x8m81  M2_M1$$202395692_3v1024x8m81_5
timestamp 1764525316
transform 1 0 680 0 1 730
box -44 -111 44 112
use M2_M1$$202395692_3v1024x8m81  M2_M1$$202395692_3v1024x8m81_6
timestamp 1764525316
transform 1 0 680 0 1 256
box -44 -111 44 112
use M2_M1$$202395692_3v1024x8m81  M2_M1$$202395692_3v1024x8m81_7
timestamp 1764525316
transform 1 0 1212 0 1 256
box -44 -111 44 112
use M2_M1$$202395692_3v1024x8m81  M2_M1$$202395692_3v1024x8m81_8
timestamp 1764525316
transform 1 0 1212 0 1 730
box -44 -111 44 112
use M2_M1$$202395692_3v1024x8m81  M2_M1$$202395692_3v1024x8m81_9
timestamp 1764525316
transform 1 0 1526 0 1 256
box -44 -111 44 112
use M2_M1$$202395692_3v1024x8m81  M2_M1$$202395692_3v1024x8m81_10
timestamp 1764525316
transform 1 0 524 0 1 1373
box -44 -111 44 112
use M2_M1$$202395692_3v1024x8m81  M2_M1$$202395692_3v1024x8m81_11
timestamp 1764525316
transform 1 0 681 0 1 1373
box -44 -111 44 112
use M2_M1$$202395692_3v1024x8m81  M2_M1$$202395692_3v1024x8m81_12
timestamp 1764525316
transform 1 0 1985 0 1 1373
box -44 -111 44 112
use M2_M1$$202395692_3v1024x8m81  M2_M1$$202395692_3v1024x8m81_13
timestamp 1764525316
transform 1 0 2613 0 1 1373
box -44 -111 44 112
use M2_M1$$202395692_3v1024x8m81  M2_M1$$202395692_3v1024x8m81_14
timestamp 1764525316
transform 1 0 1672 0 1 1373
box -44 -111 44 112
use M2_M1$$202396716_3v1024x8m81  M2_M1$$202396716_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1036 0 1 1589
box -44 -351 44 351
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2597 0 1 256
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_1
timestamp 1764525316
transform 1 0 2380 0 1 720
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_2
timestamp 1764525316
transform 1 0 2380 0 1 256
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_3
timestamp 1764525316
transform 1 0 1026 0 1 720
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_4
timestamp 1764525316
transform 1 0 1528 0 1 723
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_5
timestamp 1764525316
transform 1 0 1026 0 1 256
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_6
timestamp 1764525316
transform 1 0 0 0 1 256
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_7
timestamp 1764525316
transform 1 0 210 0 1 248
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_8
timestamp 1764525316
transform 1 0 0 0 1 720
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_9
timestamp 1764525316
transform 1 0 210 0 1 719
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_10
timestamp 1764525316
transform 1 0 0 0 1 1854
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_11
timestamp 1764525316
transform 1 0 210 0 1 1846
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_12
timestamp 1764525316
transform 1 0 210 0 1 1362
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_13
timestamp 1764525316
transform 1 0 681 0 1 1846
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_14
timestamp 1764525316
transform 1 0 0 0 1 1362
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_15
timestamp 1764525316
transform 1 0 0 0 1 1362
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_16
timestamp 1764525316
transform 1 0 2613 0 1 1876
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_17
timestamp 1764525316
transform 1 0 2299 0 1 1876
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_18
timestamp 1764525316
transform 1 0 1985 0 1 1846
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_19
timestamp 1764525316
transform 1 0 2926 0 1 1846
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_20
timestamp 1764525316
transform 1 0 3232 0 1 1362
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_21
timestamp 1764525316
transform 1 0 3294 0 1 1854
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_22
timestamp 1764525316
transform 1 0 3416 0 1 1362
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_23
timestamp 1764525316
transform 1 0 3416 0 1 1362
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_24
timestamp 1764525316
transform 1 0 2926 0 1 1332
box -45 -122 45 123
use M2_M1$$202406956_3v1024x8m81  M2_M1$$202406956_3v1024x8m81_25
timestamp 1764525316
transform 1 0 1672 0 1 1846
box -45 -122 45 123
use M2_M14310591302035_3v1024x8m81  M2_M14310591302035_3v1024x8m81_0
timestamp 1764525316
transform 1 0 520 0 1 961
box -72 -34 72 34
use M2_M14310591302035_3v1024x8m81  M2_M14310591302035_3v1024x8m81_1
timestamp 1764525316
transform 1 0 520 0 1 1122
box -72 -34 72 34
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1744 0 1 245
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_1
timestamp 1764525316
transform 1 0 2380 0 1 256
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_2
timestamp 1764525316
transform 1 0 2058 0 1 719
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_3
timestamp 1764525316
transform 1 0 2380 0 1 720
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_4
timestamp 1764525316
transform 1 0 2058 0 1 245
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_5
timestamp 1764525316
transform 1 0 2597 0 1 256
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_6
timestamp 1764525316
transform 1 0 1744 0 1 719
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_7
timestamp 1764525316
transform 1 0 1528 0 1 720
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_8
timestamp 1764525316
transform 1 0 1026 0 1 720
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_9
timestamp 1764525316
transform 1 0 0 0 1 256
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_10
timestamp 1764525316
transform 1 0 210 0 1 248
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_11
timestamp 1764525316
transform 1 0 0 0 1 720
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_12
timestamp 1764525316
transform 1 0 524 0 1 719
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_13
timestamp 1764525316
transform 1 0 680 0 1 719
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_14
timestamp 1764525316
transform 1 0 210 0 1 719
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_15
timestamp 1764525316
transform 1 0 680 0 1 245
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_16
timestamp 1764525316
transform 1 0 1212 0 1 245
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_17
timestamp 1764525316
transform 1 0 1212 0 1 719
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_18
timestamp 1764525316
transform 1 0 1526 0 1 245
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_19
timestamp 1764525316
transform 1 0 1026 0 1 256
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_20
timestamp 1764525316
transform 1 0 681 0 1 1846
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_21
timestamp 1764525316
transform 1 0 0 0 1 1854
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_22
timestamp 1764525316
transform 1 0 0 0 1 1362
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_23
timestamp 1764525316
transform 1 0 210 0 1 1846
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_24
timestamp 1764525316
transform 1 0 210 0 1 1362
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_25
timestamp 1764525316
transform 1 0 2299 0 1 1876
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_26
timestamp 1764525316
transform 1 0 1985 0 1 1846
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_27
timestamp 1764525316
transform 1 0 3232 0 1 1362
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_28
timestamp 1764525316
transform 1 0 3294 0 1 1854
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_29
timestamp 1764525316
transform 1 0 3416 0 1 1362
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_30
timestamp 1764525316
transform 1 0 2613 0 1 1876
box -45 -122 45 123
use M3_M2$$201252908_3v1024x8m81  M3_M2$$201252908_3v1024x8m81_31
timestamp 1764525316
transform 1 0 1672 0 1 1846
box -45 -122 45 123
use M3_M2$$202397740_3v1024x8m81  M3_M2$$202397740_3v1024x8m81_0
timestamp 1764525316
transform 1 0 524 0 1 1373
box -45 -112 45 112
use M3_M2$$202397740_3v1024x8m81  M3_M2$$202397740_3v1024x8m81_1
timestamp 1764525316
transform 1 0 681 0 1 1373
box -45 -112 45 112
use M3_M2$$202397740_3v1024x8m81  M3_M2$$202397740_3v1024x8m81_2
timestamp 1764525316
transform 1 0 1985 0 1 1373
box -45 -112 45 112
use M3_M2$$202397740_3v1024x8m81  M3_M2$$202397740_3v1024x8m81_3
timestamp 1764525316
transform 1 0 2613 0 1 1373
box -45 -112 45 112
use M3_M2$$202397740_3v1024x8m81  M3_M2$$202397740_3v1024x8m81_4
timestamp 1764525316
transform 1 0 1672 0 1 1373
box -45 -112 45 112
use M3_M24310591302036_3v1024x8m81  M3_M24310591302036_3v1024x8m81_0
timestamp 1764525316
transform 1 0 520 0 1 961
box -72 -35 72 35
use M3_M24310591302036_3v1024x8m81  M3_M24310591302036_3v1024x8m81_1
timestamp 1764525316
transform 1 0 520 0 1 1122
box -72 -35 72 35
use nmos_1p2$$202594348_3v1024x8m81  nmos_1p2$$202594348_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2515 0 1 1300
box -102 -44 130 171
use nmos_1p2$$202595372_3v1024x8m81  nmos_1p2$$202595372_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1417 0 1 1358
box -102 -44 130 133
use nmos_1p2$$202595372_3v1024x8m81  nmos_1p2$$202595372_3v1024x8m81_1
timestamp 1764525316
transform 1 0 1887 0 1 1358
box -102 -44 130 133
use nmos_1p2$$202596396_3v1024x8m81  nmos_1p2$$202596396_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2047 0 1 1358
box -102 -44 130 133
use nmos_1p2$$202596396_3v1024x8m81  nmos_1p2$$202596396_3v1024x8m81_1
timestamp 1764525316
transform 1 0 1577 0 1 1358
box -102 -44 130 133
use nmos_1p2$$202598444_3v1024x8m81  nmos_1p2$$202598444_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1094 0 1 1173
box -102 -44 130 255
use nmos_5p0431059130208_3v1024x8m81  nmos_5p0431059130208_3v1024x8m81_0
timestamp 1764525316
transform 1 0 419 0 -1 842
box -88 -44 144 133
use nmos_5p0431059130208_3v1024x8m81  nmos_5p0431059130208_3v1024x8m81_1
timestamp 1764525316
transform 1 0 737 0 -1 785
box -88 -44 144 133
use nmos_5p0431059130208_3v1024x8m81  nmos_5p0431059130208_3v1024x8m81_2
timestamp 1764525316
transform 1 0 259 0 -1 842
box -88 -44 144 133
use nmos_5p0431059130208_3v1024x8m81  nmos_5p0431059130208_3v1024x8m81_3
timestamp 1764525316
transform 1 0 737 0 1 1304
box -88 -44 144 133
use nmos_5p04310591302010_3v1024x8m81  nmos_5p04310591302010_3v1024x8m81_0
timestamp 1764525316
transform 1 0 3139 0 1 1173
box -88 -44 144 255
use nmos_5p04310591302039_3v1024x8m81  nmos_5p04310591302039_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2847 0 1 1173
box -116 -44 276 255
use nmos_5p04310591302040_3v1024x8m81  nmos_5p04310591302040_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1258 0 -1 785
box -88 -44 144 171
use nmos_5p04310591302040_3v1024x8m81  nmos_5p04310591302040_3v1024x8m81_1
timestamp 1764525316
transform 1 0 253 0 1 1246
box -88 -44 144 171
use nmos_5p04310591302040_3v1024x8m81  nmos_5p04310591302040_3v1024x8m81_2
timestamp 1764525316
transform 1 0 413 0 1 1246
box -88 -44 144 171
use nmos_5p04310591302042_3v1024x8m81  nmos_5p04310591302042_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1847 0 -1 785
box -144 -44 409 118
use pmos_1p2$$202583084_3v1024x8m81  pmos_1p2$$202583084_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2388 0 1 1767
box -216 -86 348 245
use pmos_1p2$$202584108_3v1024x8m81  pmos_1p2$$202584108_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1887 0 1 1687
box -188 -86 216 297
use pmos_1p2$$202585132_3v1024x8m81  pmos_1p2$$202585132_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2047 0 1 1687
box -188 -86 216 297
use pmos_1p2$$202586156_3v1024x8m81  pmos_1p2$$202586156_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1583 0 1 1687
box -188 -86 216 297
use pmos_1p2$$202587180_3v1024x8m81  pmos_1p2$$202587180_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1075 0 1 1687
box -188 -86 216 297
use pmos_5p04310591302014_3v1024x8m81  pmos_5p04310591302014_3v1024x8m81_0
timestamp 1764525316
transform 1 0 259 0 -1 401
box -174 -86 230 297
use pmos_5p04310591302014_3v1024x8m81  pmos_5p04310591302014_3v1024x8m81_1
timestamp 1764525316
transform 1 0 737 0 -1 401
box -174 -86 230 297
use pmos_5p04310591302014_3v1024x8m81  pmos_5p04310591302014_3v1024x8m81_2
timestamp 1764525316
transform 1 0 419 0 -1 401
box -174 -86 230 297
use pmos_5p04310591302014_3v1024x8m81  pmos_5p04310591302014_3v1024x8m81_3
timestamp 1764525316
transform 1 0 253 0 1 1687
box -174 -86 230 297
use pmos_5p04310591302014_3v1024x8m81  pmos_5p04310591302014_3v1024x8m81_4
timestamp 1764525316
transform 1 0 737 0 1 1687
box -174 -86 230 297
use pmos_5p04310591302014_3v1024x8m81  pmos_5p04310591302014_3v1024x8m81_5
timestamp 1764525316
transform 1 0 413 0 1 1687
box -174 -86 230 297
use pmos_5p04310591302020_3v1024x8m81  pmos_5p04310591302020_3v1024x8m81_0
timestamp 1764525316
transform 1 0 2847 0 1 1687
box -202 -86 362 297
use pmos_5p04310591302035_3v1024x8m81  pmos_5p04310591302035_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1288 0 -1 401
box -202 -86 362 245
use pmos_5p04310591302041_3v1024x8m81  pmos_5p04310591302041_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1315 0 1 1701
box -174 -86 230 175
use pmos_5p04310591302043_3v1024x8m81  pmos_5p04310591302043_3v1024x8m81_0
timestamp 1764525316
transform 1 0 1850 0 -1 401
box -230 -86 495 272
<< labels >>
rlabel metal3 s 95 743 95 743 4 vss
port 1 nsew
rlabel metal3 s 454 956 454 956 4 GWEN
port 2 nsew
rlabel metal3 s 95 1362 95 1362 4 vss
port 1 nsew
rlabel metal3 s 95 1846 95 1846 4 vdd
port 3 nsew
rlabel metal3 s 454 1117 454 1117 4 VSS
port 4 nsew
rlabel metal3 s 95 301 95 301 4 vdd
port 3 nsew
rlabel metal1 s 249 2162 249 2162 4 men
port 5 nsew
rlabel metal1 s 2215 560 2215 560 4 wep
port 6 nsew
rlabel metal1 s 101 21 101 21 4 wen
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 3403 2300
string MASKHINTS_PPLUS 133 1641 3155 1974 139 144 913 447 1139 169 2291 448
string path 15.820 2.690 15.820 4.995 
<< end >>
