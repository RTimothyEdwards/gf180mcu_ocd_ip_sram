magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nwell >>
rect -133 -66 160 1039
<< polysilicon >>
rect -14 973 41 1007
rect -14 -34 41 0
use pmos_5p04310591302072_3v256x8m81  pmos_5p04310591302072_3v256x8m81_0
timestamp 1763766357
transform 1 0 -14 0 1 0
box -174 -86 230 1059
<< end >>
