magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< nwell >>
rect -41 8409 610 11860
rect -13 4936 627 5174
rect -130 4924 627 4936
rect -130 4481 609 4924
rect -48 4479 609 4481
<< pmos >>
rect 172 10921 228 11239
rect 332 10921 388 11239
rect 172 10416 228 10733
rect 332 10416 388 10733
rect 67 4568 123 4707
rect 319 4568 375 4707
<< pdiff >>
rect 46 11195 172 11239
rect 46 11149 97 11195
rect 143 11149 172 11195
rect 46 11013 172 11149
rect 46 10967 97 11013
rect 143 10967 172 11013
rect 46 10921 172 10967
rect 228 11195 332 11239
rect 228 11149 257 11195
rect 303 11149 332 11195
rect 228 11013 332 11149
rect 228 10967 257 11013
rect 303 10967 332 11013
rect 228 10921 332 10967
rect 388 11195 523 11239
rect 388 11149 443 11195
rect 489 11149 523 11195
rect 388 11013 523 11149
rect 388 10967 443 11013
rect 489 10967 523 11013
rect 388 10921 523 10967
rect 46 10690 172 10733
rect 46 10644 97 10690
rect 143 10644 172 10690
rect 46 10508 172 10644
rect 46 10462 97 10508
rect 143 10462 172 10508
rect 46 10416 172 10462
rect 228 10690 332 10733
rect 228 10644 257 10690
rect 303 10644 332 10690
rect 228 10508 332 10644
rect 228 10462 257 10508
rect 303 10462 332 10508
rect 228 10416 332 10462
rect 388 10690 523 10733
rect 388 10644 443 10690
rect 489 10644 523 10690
rect 388 10508 523 10644
rect 388 10462 443 10508
rect 489 10462 523 10508
rect 388 10416 523 10462
rect -44 4662 67 4707
rect -44 4615 -24 4662
rect 22 4615 67 4662
rect -44 4568 67 4615
rect 123 4661 319 4707
rect 123 4615 208 4661
rect 254 4615 319 4661
rect 123 4568 319 4615
rect 375 4661 523 4707
rect 375 4615 447 4661
rect 493 4615 523 4661
rect 375 4568 523 4615
<< pdiffc >>
rect 97 11149 143 11195
rect 97 10967 143 11013
rect 257 11149 303 11195
rect 257 10967 303 11013
rect 443 11149 489 11195
rect 443 10967 489 11013
rect 97 10644 143 10690
rect 97 10462 143 10508
rect 257 10644 303 10690
rect 257 10462 303 10508
rect 443 10644 489 10690
rect 443 10462 489 10508
rect -24 4615 22 4662
rect 208 4615 254 4661
rect 447 4615 493 4661
<< nsubdiff >>
rect 119 11552 523 11712
<< polysilicon >>
rect 172 11239 228 11436
rect 332 11239 388 11436
rect 172 10733 228 10921
rect 332 10733 388 10921
rect 172 10352 228 10416
rect 332 10352 388 10416
rect 172 10268 388 10352
rect 218 10267 304 10268
rect 248 10119 304 10267
rect 250 8475 306 8555
rect 250 6866 306 7513
rect 250 6045 306 6152
rect 250 5851 306 5952
rect 67 4848 375 4947
rect 67 4707 123 4848
rect 319 4707 375 4848
rect 67 4543 123 4568
rect 67 4470 194 4543
rect 319 4532 375 4568
rect 138 4410 194 4470
rect 306 4470 375 4532
rect 306 4410 362 4470
rect 138 4243 194 4272
rect 306 4243 362 4272
<< metal1 >>
rect 49 11562 523 11717
rect 74 11434 494 11562
rect 74 11195 159 11434
rect 74 11149 97 11195
rect 143 11149 159 11195
rect 74 11013 159 11149
rect 74 10967 97 11013
rect 143 10967 159 11013
rect 74 10690 159 10967
rect 222 11195 337 11382
rect 222 11149 257 11195
rect 303 11149 337 11195
rect 222 11013 337 11149
rect 222 10967 257 11013
rect 303 10967 337 11013
rect 222 10930 337 10967
rect 402 11195 494 11434
rect 402 11149 443 11195
rect 489 11149 494 11195
rect 402 11013 494 11149
rect 402 10967 443 11013
rect 489 10967 494 11013
rect 74 10644 97 10690
rect 143 10644 159 10690
rect 74 10508 159 10644
rect 74 10462 97 10508
rect 143 10462 159 10508
rect 74 10425 159 10462
rect 222 10690 337 10879
rect 222 10644 257 10690
rect 303 10644 337 10690
rect 222 10508 337 10644
rect 222 10462 257 10508
rect 303 10462 337 10508
rect 222 10425 337 10462
rect 402 10690 494 10967
rect 402 10644 443 10690
rect 489 10644 494 10690
rect 402 10508 494 10644
rect 402 10462 443 10508
rect 489 10462 494 10508
rect 402 10425 494 10462
rect 68 9710 219 9890
rect 333 9710 494 9890
rect 119 9065 182 9231
rect 130 8751 182 9065
rect 119 8647 182 8751
rect 119 7557 189 8647
rect 236 8296 332 8479
rect 381 7497 445 9227
rect 45 7381 445 7497
rect 43 7103 523 7237
rect 113 6958 379 7055
rect 113 6191 188 6958
rect 380 6232 457 6816
rect 113 5187 181 6191
rect 239 6031 331 6124
rect 239 5873 331 5966
rect 378 5193 457 6232
rect -41 5001 73 5085
rect -41 4662 31 5001
rect 198 4858 374 4955
rect -41 4615 -24 4662
rect 22 4615 31 4662
rect -41 4577 31 4615
rect 205 4661 288 4777
rect 205 4615 208 4661
rect 254 4615 288 4661
rect 37 4218 120 4433
rect 205 4313 288 4615
rect 443 4661 523 5085
rect 443 4615 447 4661
rect 493 4615 523 4661
rect 443 4577 523 4615
rect 378 4218 457 4433
rect 37 4096 457 4218
<< metal2 >>
rect 68 11314 124 11715
rect 216 11435 344 11717
rect 245 11434 344 11435
rect 68 11258 327 11314
rect 68 9109 124 11258
rect 438 10808 494 11715
rect 285 10752 494 10808
rect 248 7368 304 8406
rect 143 7312 304 7368
rect 143 5938 199 7312
rect 438 7073 494 10752
rect 256 7013 494 7073
rect 411 6124 474 6956
rect 260 6027 474 6124
rect 143 5882 312 5938
rect 143 4777 199 5882
rect 411 5494 474 6027
rect 270 5397 474 5494
rect 270 4858 330 5397
rect 143 4597 290 4777
rect 172 4063 272 4211
<< metal3 >>
rect -65 10338 525 11716
rect -41 7127 525 8527
rect -41 6881 525 7021
rect -41 6639 525 6779
rect -41 6398 525 6538
rect -41 6156 525 6296
rect -41 5924 525 6064
rect -41 5682 525 5822
rect -41 5440 525 5580
rect -41 5198 525 5338
rect -41 4610 525 5052
rect -41 4017 525 4464
use M1_NWELL05_512x8m81  M1_NWELL05_512x8m81_0
timestamp 1763564386
transform 1 0 285 0 1 11632
box -265 -159 265 159
use M1_NWELL09_512x8m81  M1_NWELL09_512x8m81_1
timestamp 1763564386
transform 1 0 279 0 1 5043
box -320 -159 320 159
use M1_POLY24310591302030_512x8m81  M1_POLY24310591302030_512x8m81_0
timestamp 1763564386
transform 1 0 272 0 1 10310
box -95 -36 95 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1763564386
transform 1 0 253 0 1 4905
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1763564386
transform 1 0 290 0 1 5910
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_2
timestamp 1763564386
transform 1 0 281 0 1 6087
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_6
timestamp 1763564386
transform 1 0 276 0 1 8442
box -36 -36 36 36
use M1_PSUB$$45111340_512x8m81  M1_PSUB$$45111340_512x8m81_0
timestamp 1763564386
transform 1 0 120 0 1 7168
box -56 -58 56 58
use M1_PSUB$$45111340_512x8m81  M1_PSUB$$45111340_512x8m81_1
timestamp 1763564386
transform 1 0 435 0 1 7168
box -56 -58 56 58
use M1_PSUB$$47122476_512x8m81  M1_PSUB$$47122476_512x8m81_0
timestamp 1763564386
transform 1 0 269 0 1 4160
box -223 -58 254 57
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_0
timestamp 1763564386
transform 1 0 247 0 1 4689
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_2
timestamp 1763564386
transform 1 0 106 0 1 9800
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_3
timestamp 1763564386
transform 1 0 108 0 1 9168
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_4
timestamp 1763564386
transform 1 0 281 0 1 11285
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_5
timestamp 1763564386
transform 1 0 276 0 1 8389
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_6
timestamp 1763564386
transform 1 0 456 0 1 9800
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_7
timestamp 1763564386
transform 1 0 281 0 1 10780
box -34 -63 34 63
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_0
timestamp 1763564386
transform 1 0 304 0 1 4904
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_1
timestamp 1763564386
transform 1 0 295 0 1 5910
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_5
timestamp 1763564386
transform 0 1 117 -1 0 7460
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_6
timestamp 1763564386
transform 1 0 344 0 1 7185
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_9
timestamp 1763564386
transform 1 0 291 0 1 6994
box -35 -56 35 55
use M3_M2431059130201_512x8m81  M3_M2431059130201_512x8m81_1
timestamp 1763564386
transform 1 0 344 0 1 7192
box -35 -63 35 63
use nmos_1p2$$47119404_512x8m81  nmos_1p2$$47119404_512x8m81_1
timestamp 1763564386
transform 1 0 264 0 -1 6826
box -102 -44 130 679
use nmos_1p2$$47119404_512x8m81  nmos_1p2$$47119404_512x8m81_3
timestamp 1763564386
transform 1 0 264 0 -1 8190
box -102 -44 130 679
use nmos_5p0431059130202_512x8m81  nmos_5p0431059130202_512x8m81_0
timestamp 1763564386
transform 1 0 170 0 1 4315
box -124 -44 285 98
use pmos_1p2$$46889004_512x8m81  pmos_1p2$$46889004_512x8m81_1
timestamp 1763564386
transform 1 0 264 0 -1 5811
box -188 -86 216 721
use pmos_5p0431059130201_512x8m81  pmos_5p0431059130201_512x8m81_0
timestamp 1763564386
transform 1 0 248 0 -1 10077
box -174 -86 230 721
use pmos_5p0431059130201_512x8m81  pmos_5p0431059130201_512x8m81_1
timestamp 1763564386
transform 1 0 250 0 -1 9231
box -174 -86 230 721
use via1_2_512x8m81  via1_2_512x8m81_0
timestamp 1763564386
transform 1 0 174 0 1 4115
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_0
timestamp 1763564386
transform 1 0 259 0 1 6029
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_2
timestamp 1763564386
transform 0 -1 343 1 0 11435
box 0 0 65 89
use via1_R90_512x8m81  via1_R90_512x8m81_3
timestamp 1763564386
transform 0 -1 343 1 0 11621
box 0 0 65 89
use via2_R90_512x8m81  via2_R90_512x8m81_0
timestamp 1763564386
transform 0 -1 373 1 0 11435
box 0 0 65 89
use via2_R90_512x8m81  via2_R90_512x8m81_1
timestamp 1763564386
transform 0 -1 373 1 0 11621
box 0 0 65 89
<< labels >>
rlabel metal1 s 229 10312 229 10312 4 pcb
port 8 nsew
rlabel metal2 s 105 11421 105 11421 4 bb
port 4 nsew
rlabel metal2 s 428 11421 428 11421 4 b
port 3 nsew
rlabel metal3 s 318 11384 318 11384 4 vdd
port 2 nsew
rlabel metal2 s 281 4925 281 4925 4 ypass
port 6 nsew
rlabel metal1 s 318 5059 318 5059 4 vdd
port 2 nsew
rlabel metal3 s 303 6426 303 6426 4 vss
port 1 nsew
<< properties >>
string path 0.000 27.385 0.000 -0.005 
<< end >>
