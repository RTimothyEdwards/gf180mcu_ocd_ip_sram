magic
tech gf180mcuD
magscale 1 5
timestamp 1763765945
<< metal1 >>
rect -133 13 133 23
rect -133 -13 -124 13
rect 124 -13 133 13
rect -133 -23 133 -13
<< via1 >>
rect -124 -13 124 13
<< metal2 >>
rect -133 13 133 23
rect -133 -13 -124 13
rect 124 -13 133 13
rect -133 -23 133 -13
<< end >>
