magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal1 >>
rect -44 731 38 732
rect -44 711 44 731
rect -44 -711 -26 711
rect 26 -711 44 711
rect -44 -732 44 -711
<< via1 >>
rect -26 -711 26 711
<< metal2 >>
rect -44 711 44 731
rect -44 -711 -26 711
rect 26 -711 44 711
rect -44 -732 44 -711
<< end >>
