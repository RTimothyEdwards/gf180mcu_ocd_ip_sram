magic
tech gf180mcuD
magscale 1 10
timestamp 1763657283
<< metal2 >>
rect 20083 4542 20393 4960
rect 41878 4584 42188 4915
use M2_M14310591302012_256x8m81  M2_M14310591302012_256x8m81_0
timestamp 1763564386
transform 1 0 42036 0 1 4752
box -113 -156 113 156
use M2_M14310591302012_256x8m81  M2_M14310591302012_256x8m81_1
timestamp 1763564386
transform 1 0 20240 0 1 4752
box -113 -156 113 156
use M3_M2431059130206_256x8m81  M3_M2431059130206_256x8m81_0
timestamp 1763564386
transform 1 0 42036 0 1 4751
box -113 -156 113 156
use M3_M2431059130206_256x8m81  M3_M2431059130206_256x8m81_1
timestamp 1763564386
transform 1 0 20240 0 1 4711
box -113 -156 113 156
use power_route_01_256x8m81  power_route_01_256x8m81_0
timestamp 1763564386
transform -1 0 59708 0 1 46637
box -357 0 1199 1697
use power_route_01_256x8m81  power_route_01_256x8m81_1
timestamp 1763564386
transform -1 0 18635 0 1 46637
box -357 0 1199 1697
use power_route_01_256x8m81  power_route_01_256x8m81_2
timestamp 1763564386
transform 1 0 6623 0 1 46637
box -357 0 1199 1697
use power_route_01_256x8m81  power_route_01_256x8m81_3
timestamp 1763564386
transform 1 0 14443 0 1 46637
box -357 0 1199 1697
use power_route_01_256x8m81  power_route_01_256x8m81_4
timestamp 1763564386
transform 1 0 10533 0 1 46637
box -357 0 1199 1697
use power_route_01_256x8m81  power_route_01_256x8m81_5
timestamp 1763564386
transform 1 0 43806 0 1 46637
box -357 0 1199 1697
use power_route_01_256x8m81  power_route_01_256x8m81_6
timestamp 1763564386
transform 1 0 55526 0 1 46637
box -357 0 1199 1697
use power_route_01_256x8m81  power_route_01_256x8m81_7
timestamp 1763564386
transform 1 0 51616 0 1 46637
box -357 0 1199 1697
use power_route_01_256x8m81  power_route_01_256x8m81_8
timestamp 1763564386
transform 1 0 47714 0 1 46637
box -357 0 1199 1697
use power_route_01_256x8m81  power_route_01_256x8m81_9
timestamp 1763564386
transform 1 0 2713 0 1 46637
box -357 0 1199 1697
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_15
timestamp 1763564386
transform 1 0 -992 0 1 46054
box 2337 -175 21427 945
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_16
timestamp 1763564386
transform 1 0 -992 0 1 44842
box 2337 -175 21427 945
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_17
timestamp 1763564386
transform 1 0 -992 0 1 42418
box 2337 -175 21427 945
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_18
timestamp 1763564386
transform 1 0 -992 0 1 43630
box 2337 -175 21427 945
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_19
timestamp 1763564386
transform 1 0 -992 0 1 37570
box 2337 -175 21427 945
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_20
timestamp 1763564386
transform 1 0 -992 0 1 38782
box 2337 -175 21427 945
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_21
timestamp 1763564386
transform 1 0 -992 0 1 41206
box 2337 -175 21427 945
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_22
timestamp 1763564386
transform 1 0 -992 0 1 39994
box 2337 -175 21427 945
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_23
timestamp 1763564386
transform 1 0 -992 0 1 36358
box 2337 -175 21427 945
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_24
timestamp 1763564386
transform 1 0 -992 0 1 35146
box 2337 -175 21427 945
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_25
timestamp 1763564386
transform 1 0 -992 0 1 32722
box 2337 -175 21427 945
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_26
timestamp 1763564386
transform 1 0 -992 0 1 33934
box 2337 -175 21427 945
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_27
timestamp 1763564386
transform 1 0 -992 0 1 27874
box 2337 -175 21427 945
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_28
timestamp 1763564386
transform 1 0 -992 0 1 29086
box 2337 -175 21427 945
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_29
timestamp 1763564386
transform 1 0 -992 0 1 31510
box 2337 -175 21427 945
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_30
timestamp 1763564386
transform 1 0 -992 0 1 30298
box 2337 -175 21427 945
use power_route_02_a_256x8m81  power_route_02_a_256x8m81_31
timestamp 1763564386
transform 1 0 -992 0 1 26662
box 2337 -175 21427 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_0
timestamp 1763565237
transform -1 0 64142 0 1 27871
box 2538 -155 21443 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_1
timestamp 1763565237
transform -1 0 64142 0 1 29083
box 2538 -155 21443 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_2
timestamp 1763565237
transform -1 0 64142 0 1 30295
box 2538 -155 21443 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_3
timestamp 1763565237
transform -1 0 64142 0 1 31507
box 2538 -155 21443 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_4
timestamp 1763565237
transform -1 0 64142 0 1 32719
box 2538 -155 21443 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_5
timestamp 1763565237
transform -1 0 64142 0 1 33931
box 2538 -155 21443 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_6
timestamp 1763565237
transform -1 0 64142 0 1 35143
box 2538 -155 21443 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_7
timestamp 1763565237
transform -1 0 64142 0 1 36355
box 2538 -155 21443 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_8
timestamp 1763565237
transform -1 0 64142 0 1 37567
box 2538 -155 21443 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_9
timestamp 1763565237
transform -1 0 64142 0 1 38779
box 2538 -155 21443 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_10
timestamp 1763565237
transform -1 0 64142 0 1 39991
box 2538 -155 21443 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_11
timestamp 1763565237
transform -1 0 64142 0 1 41203
box 2538 -155 21443 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_12
timestamp 1763565237
transform -1 0 64142 0 1 42415
box 2538 -155 21443 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_13
timestamp 1763565237
transform -1 0 64142 0 1 43627
box 2538 -155 21443 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_14
timestamp 1763565237
transform -1 0 64142 0 1 44839
box 2538 -155 21443 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_15
timestamp 1763565237
transform -1 0 64142 0 1 46051
box 2538 -155 21443 945
use power_route_02_b_256x8m81  power_route_02_b_256x8m81_32
timestamp 1763565237
transform -1 0 64142 0 1 26659
box 2538 -155 21443 945
use power_route_04_256x8m81  power_route_04_256x8m81_0
timestamp 1763578215
transform -1 0 63942 0 1 170
box 2338 4041 4642 36851
use power_route_04_256x8m81  power_route_04_256x8m81_1
timestamp 1763578215
transform 1 0 -992 0 1 170
box 2338 4041 4642 36851
use power_route_05_256x8m81  power_route_05_256x8m81_0
timestamp 1763564386
transform 1 0 14119 0 1 1725
box -5 1821 864 5538
use power_route_05_256x8m81  power_route_05_256x8m81_1
timestamp 1763564386
transform 1 0 47412 0 1 1725
box -5 1821 864 5538
use power_route_05_256x8m81  power_route_05_256x8m81_2
timestamp 1763564386
transform 1 0 55242 0 1 1721
box -5 1821 864 5538
use power_route_05_256x8m81  power_route_05_256x8m81_3
timestamp 1763564386
transform 1 0 6357 0 1 1725
box -5 1821 864 5538
use power_route_06_256x8m81  power_route_06_256x8m81_0
timestamp 1763578215
transform 1 0 42568 0 1 1321
box -4 2229 863 13188
use power_route_06_256x8m81  power_route_06_256x8m81_1
timestamp 1763578215
transform 1 0 18748 0 1 1315
box -4 2229 863 13188
use power_route_07_256x8m81  power_route_07_256x8m81_0
timestamp 1763580222
transform 1 0 28522 0 1 1725
box -5 2486 864 4904
use power_route_07_256x8m81  power_route_07_256x8m81_1
timestamp 1763580222
transform 1 0 27248 0 1 1725
box -5 2486 864 4904
<< end >>
