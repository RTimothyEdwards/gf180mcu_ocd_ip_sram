magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal1 >>
rect -1782 156 1782 165
rect -1782 -156 -1773 156
rect 1773 -156 1782 156
rect -1782 -165 1782 -156
<< via1 >>
rect -1773 -156 1773 156
<< metal2 >>
rect -1782 156 1782 165
rect -1782 -156 -1773 156
rect 1773 -156 1782 156
rect -1782 -165 1782 -156
<< end >>
