magic
tech gf180mcuD
magscale 1 10
timestamp 1763575302
<< metal2 >>
rect -113 1148 113 1155
rect -113 -648 -106 1148
rect 106 -648 113 1148
rect -113 -655 113 -648
<< via2 >>
rect -106 -648 106 1148
<< metal3 >>
rect -113 1148 113 1155
rect -113 -648 -106 1148
rect 106 -648 113 1148
rect -113 -655 113 -648
<< end >>
