magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< nwell >>
rect -133 -65 160 1124
<< polysilicon >>
rect -14 1058 41 1087
rect -14 -34 41 0
use pmos_5p04310591302068_3v1024x8m81  pmos_5p04310591302068_3v1024x8m81_0
timestamp 1764525316
transform 1 0 -14 0 1 0
box -174 -86 230 1144
<< end >>
