magic
tech gf180mcuD
magscale 1 10
timestamp 1763570009
<< nwell >>
rect -100 -1819 774 -1500
<< nmos >>
rect 145 -4624 201 -3988
rect 305 -4624 361 -3988
rect 465 -4624 521 -3988
<< ndiff >>
rect 54 -4001 145 -3988
rect 54 -4564 70 -4001
rect 116 -4564 145 -4001
rect 54 -4624 145 -4564
rect 201 -4624 305 -3988
rect 361 -4624 465 -3988
rect 521 -4001 618 -3988
rect 521 -4564 550 -4001
rect 597 -4564 618 -4001
rect 521 -4624 618 -4564
<< ndiffc >>
rect 70 -4564 116 -4001
rect 550 -4564 597 -4001
<< psubdiff >>
rect 0 138 674 171
rect 0 91 141 138
rect 520 91 674 138
rect 0 56 674 91
rect 0 -4810 674 -4776
rect 0 -4857 141 -4810
rect 519 -4857 674 -4810
rect 0 -4891 674 -4857
<< nsubdiff >>
rect 0 -1637 674 -1604
rect 0 -1683 133 -1637
rect 401 -1683 674 -1637
rect 0 -1716 674 -1683
<< psubdiffcont >>
rect 141 91 520 138
rect 141 -4857 519 -4810
<< nsubdiffcont >>
rect 133 -1683 401 -1637
<< polysilicon >>
rect 145 -475 201 -342
rect 305 -475 361 -342
rect 465 -475 521 -342
rect 145 -539 521 -475
rect 145 -566 201 -539
rect 305 -566 361 -539
rect 465 -566 521 -539
rect 145 -1459 201 -1184
rect 305 -1459 361 -1184
rect 465 -1459 521 -1184
rect 145 -1517 521 -1459
rect 145 -3988 201 -2751
rect 305 -3988 361 -2751
rect 465 -3988 521 -2751
rect 145 -4683 201 -4624
rect 305 -4683 361 -4624
rect 465 -4683 521 -4624
<< metal1 >>
rect 0 138 674 165
rect 0 91 141 138
rect 520 91 674 138
rect 0 -38 674 91
rect 60 -175 142 -38
rect 374 -175 455 -38
rect 217 -465 298 -354
rect 217 -466 301 -465
rect 531 -466 611 -230
rect 217 -499 611 -466
rect 218 -549 611 -499
rect 218 -651 298 -549
rect 531 -651 611 -549
rect 140 -1536 611 -1453
rect 0 -1637 455 -1618
rect 0 -1683 133 -1637
rect 401 -1683 455 -1637
rect 0 -1701 455 -1683
rect 60 -1913 142 -1701
rect 374 -1914 455 -1701
rect 531 -2254 611 -1536
rect -40 -2861 714 -2797
rect -40 -3003 714 -2938
rect -40 -3144 714 -3080
rect -40 -3285 714 -3221
rect -40 -3426 714 -3362
rect -40 -3567 714 -3503
rect 60 -4001 142 -3973
rect 60 -4564 70 -4001
rect 116 -4564 142 -4001
rect 60 -4680 142 -4564
rect 531 -4001 612 -3973
rect 531 -4564 550 -4001
rect 597 -4485 612 -4001
rect 597 -4564 611 -4485
rect 531 -4618 611 -4564
rect 5 -4810 674 -4680
rect 5 -4857 141 -4810
rect 519 -4857 674 -4810
rect 5 -4885 674 -4857
<< metal2 >>
rect 212 -257 301 228
rect 213 -2704 616 -2459
rect 526 -2705 616 -2704
rect 527 -3882 616 -2705
<< metal3 >>
rect -36 -436 774 228
rect -40 -2727 757 -908
rect 0 -4986 674 -3700
use M1_POLY24310591302030_256x8m81  M1_POLY24310591302030_256x8m81_0
timestamp 1763564386
transform 1 0 346 0 1 -1495
box -95 -36 95 36
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_0
timestamp 1763564386
transform 1 0 258 0 1 -2581
box -43 -122 43 122
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_1
timestamp 1763564386
transform 1 0 571 0 1 -2581
box -43 -122 43 122
use M2_M1$$43378732_256x8m81  M2_M1$$43378732_256x8m81_0
timestamp 1763564386
transform 1 0 412 0 1 -2036
box -44 -351 44 351
use M2_M1$$43378732_256x8m81  M2_M1$$43378732_256x8m81_1
timestamp 1763564386
transform 1 0 571 0 1 -4134
box -44 -351 44 351
use M2_M1$$43379756_256x8m81  M2_M1$$43379756_256x8m81_0
timestamp 1763564386
transform 1 0 415 0 1 -130
box -44 -275 44 275
use M2_M1$$43379756_256x8m81  M2_M1$$43379756_256x8m81_1
timestamp 1763564386
transform 1 0 93 0 1 -130
box -44 -275 44 275
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_0
timestamp 1763570009
transform 1 0 256 0 1 -299
box -44 -198 44 198
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_1
timestamp 1763570009
transform 1 0 415 0 1 -1107
box -44 -198 44 198
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_2
timestamp 1763570009
transform 1 0 93 0 1 -1107
box -44 -198 44 198
use M2_M1$$47515692_256x8m81  M2_M1$$47515692_256x8m81_0
timestamp 1763564386
transform 1 0 93 0 1 -2188
box -44 -504 44 284
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_0
timestamp 1763564386
transform 1 0 415 0 1 -1107
box -45 -198 45 198
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_1
timestamp 1763564386
transform 1 0 93 0 1 -1107
box -45 -198 45 198
use M3_M2$$47332396_256x8m81  M3_M2$$47332396_256x8m81_0
timestamp 1763564386
transform 1 0 93 0 1 -2188
box -45 -504 45 504
use M3_M2$$47333420_256x8m81  M3_M2$$47333420_256x8m81_0
timestamp 1763564386
transform 1 0 93 0 1 -130
box -84 -185 84 275
use M3_M2$$47333420_256x8m81  M3_M2$$47333420_256x8m81_1
timestamp 1763564386
transform 1 0 415 0 1 -130
box -84 -185 84 275
use M3_M2$$47819820_256x8m81  M3_M2$$47819820_256x8m81_0
timestamp 1763564386
transform 1 0 412 0 1 -2036
box -45 -351 45 351
use nmos_1p2$$46551084_256x8m81  nmos_1p2$$46551084_256x8m81_0
timestamp 1763564386
transform -1 0 187 0 -1 -95
box -102 -44 130 255
use nmos_1p2$$46551084_256x8m81  nmos_1p2$$46551084_256x8m81_1
timestamp 1763564386
transform -1 0 347 0 -1 -95
box -102 -44 130 255
use nmos_1p2$$46551084_256x8m81  nmos_1p2$$46551084_256x8m81_2
timestamp 1763564386
transform 1 0 479 0 -1 -95
box -102 -44 130 255
use pmos_1p2$$47820844_256x8m81  pmos_1p2$$47820844_256x8m81_0
timestamp 1763564386
transform 1 0 479 0 -1 -609
box -188 -86 216 624
use pmos_1p2$$47820844_256x8m81  pmos_1p2$$47820844_256x8m81_1
timestamp 1763564386
transform -1 0 187 0 -1 -609
box -188 -86 216 624
use pmos_1p2$$47820844_256x8m81  pmos_1p2$$47820844_256x8m81_2
timestamp 1763564386
transform -1 0 347 0 -1 -609
box -188 -86 216 624
use pmos_1p2$$47821868_256x8m81  pmos_1p2$$47821868_256x8m81_0
timestamp 1763564386
transform 1 0 159 0 1 -2710
box -188 -86 216 615
use pmos_1p2$$47821868_256x8m81  pmos_1p2$$47821868_256x8m81_2
timestamp 1763564386
transform 1 0 319 0 1 -2710
box -188 -86 216 615
use pmos_1p2$$47821868_256x8m81  pmos_1p2$$47821868_256x8m81_3
timestamp 1763564386
transform 1 0 479 0 1 -2710
box -188 -86 216 615
<< end >>
