magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< metal2 >>
rect -45 28 783 46
rect -45 -28 -28 28
rect 766 -28 783 28
rect -45 -46 783 -28
<< via2 >>
rect -28 -28 766 28
<< metal3 >>
rect -45 28 783 46
rect -45 -28 -28 28
rect 766 -28 783 28
rect -45 -46 783 -28
<< end >>
