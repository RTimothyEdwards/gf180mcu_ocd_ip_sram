magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< polysilicon >>
rect -14 615 41 648
rect -14 -33 41 0
use nmos_5p043105913020102_3v512x8m81  nmos_5p043105913020102_3v512x8m81_0
timestamp 1764525316
transform 1 0 -14 0 1 0
box -88 -44 144 659
<< end >>
