magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< error_s >>
rect 15698 -9996 15855 -9824
rect 15870 -10314 15990 -9996
<< nwell >>
rect 15513 -2147 15942 -674
rect 15513 -4026 16041 -2147
rect 15684 -6739 16071 -6535
rect 15684 -7092 16041 -6739
rect 15684 -7172 16040 -7092
rect 15713 -7951 16040 -7172
rect 15855 -9996 16474 -9613
rect 15855 -10314 15870 -9996
rect 16400 -10314 16474 -9996
rect 15855 -10335 16474 -10314
rect 15876 -10336 16474 -10335
rect 15880 -13577 15896 -13176
rect 15880 -13729 16460 -13577
rect 15879 -14859 16170 -14540
<< polysilicon >>
rect -535 39998 -439 40070
rect -535 38962 -439 39034
rect -535 38786 -439 38858
rect -535 37750 -439 37822
rect -535 37574 -439 37646
rect -535 36538 -439 36610
rect -535 36362 -439 36434
rect -535 35326 -439 35398
rect -535 35150 -439 35222
rect -535 34114 -439 34186
rect -535 33938 -439 34010
rect -535 32902 -439 32974
rect -535 32726 -439 32798
rect -535 31690 -439 31762
rect -535 31514 -439 31586
rect -535 30478 -439 30550
rect -535 30302 -439 30374
rect -535 29266 -439 29338
rect -535 29090 -439 29162
rect -535 28054 -439 28126
rect -535 27878 -439 27950
rect -535 26842 -439 26914
rect -535 26666 -439 26738
rect -535 25630 -439 25702
rect -535 25454 -439 25526
rect -535 24418 -439 24490
rect -535 24242 -439 24314
rect -535 23206 -439 23278
rect -535 23030 -439 23102
rect -535 21994 -439 22066
rect -535 21818 -439 21890
rect -535 20782 -439 20854
rect -535 20606 -439 20678
rect -535 19570 -439 19642
rect -535 19394 -439 19466
rect -535 18358 -439 18430
rect -535 18182 -439 18254
rect -535 17146 -439 17218
rect -535 16970 -439 17042
rect -535 15934 -439 16006
rect -535 15758 -439 15830
rect -535 14722 -439 14794
rect -535 14546 -439 14618
rect -535 13510 -439 13582
rect -535 13334 -439 13406
rect -535 12298 -439 12370
rect -535 12122 -439 12194
rect -535 11086 -439 11158
rect -535 10910 -439 10982
rect -535 9874 -439 9946
rect -535 9698 -439 9770
rect -535 8662 -439 8734
rect -535 8486 -439 8558
rect -535 7450 -439 7522
rect -535 7274 -439 7346
rect -535 6238 -439 6310
rect -535 6062 -439 6134
rect -535 5026 -439 5098
rect -535 4850 -439 4922
rect -535 3814 -439 3886
rect -535 3638 -439 3710
rect -535 2602 -439 2674
rect -535 2426 -439 2498
rect -535 1390 -439 1462
rect -535 1214 -439 1286
rect -535 178 -439 250
rect 16067 -10288 16123 -10269
rect 16227 -10288 16283 -10269
rect 16067 -10384 16283 -10288
rect 16067 -10481 16123 -10384
rect 16227 -10481 16283 -10384
rect 16070 -12352 16126 -12332
rect 16230 -12352 16286 -12332
rect 16070 -12444 16286 -12352
rect 16070 -12468 16126 -12444
rect 16230 -12468 16286 -12444
<< metal1 >>
rect 16572 35210 16609 35350
rect 16624 35210 16894 35350
rect -525 -240 -472 80
rect -525 -320 -275 -240
rect 16172 -3925 16353 -3213
rect 15820 -7281 16217 -7197
rect 15820 -8454 15901 -7281
rect 16357 -7557 16527 -7349
rect 15820 -8538 16522 -8454
rect 16134 -10286 16216 -10016
rect 15853 -10338 16216 -10286
rect 16440 -10296 16522 -8538
rect 15853 -12380 15904 -10338
rect 16134 -10587 16216 -10338
rect 16285 -10380 16522 -10296
rect 15977 -12257 16059 -10608
rect 16291 -12257 16373 -10608
rect 15977 -12380 16059 -12379
rect 15853 -12432 16062 -12380
rect 15981 -14741 16062 -13403
rect 16137 -13801 16219 -12830
rect 16294 -14676 16375 -13422
rect 16294 -14722 16299 -14676
rect 16345 -14722 16375 -14676
rect 16294 -14741 16375 -14722
rect 16100 -16182 16256 -14859
<< metal2 >>
rect -528 93 -472 40214
rect 16574 38797 16661 40245
rect 16123 -599 16207 113
rect 16076 -668 16207 -599
rect 16333 -599 16417 112
rect 16574 21 16661 37818
rect 16333 -668 16422 -599
rect 16076 -795 16132 -668
rect 16366 -795 16422 -668
rect 16134 -16314 16225 -12238
<< metal3 >>
rect -631 83 -432 180
rect 15604 -1898 16729 -718
rect 15446 -1957 16729 -1898
rect 15446 -2095 16727 -1957
rect 15668 -5306 16729 -3922
rect 15667 -5552 16729 -5402
rect 15667 -5798 16729 -5647
rect 15667 -6043 16729 -5892
rect 15667 -6288 16729 -6137
rect 15667 -6510 16507 -6360
rect 15667 -6752 16507 -6601
rect 15667 -7002 16507 -6852
rect 15667 -7247 16507 -7095
rect 15668 -7702 16507 -7393
rect 15604 -8416 16584 -8101
rect 15668 -8420 16584 -8416
rect 15698 -11027 16382 -9120
rect 15698 -13079 16382 -11227
rect 15698 -13549 16382 -13209
rect 15645 -13711 16382 -13549
rect 15645 -14640 16382 -14072
rect 15698 -15942 16135 -15021
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_0
timestamp 1763765945
transform -1 0 99 0 1 7836
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1
timestamp 1763765945
transform -1 0 99 0 1 2988
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_2
timestamp 1763765945
transform -1 0 99 0 1 5412
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_3
timestamp 1763765945
transform -1 0 99 0 1 10260
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_4
timestamp 1763765945
transform -1 0 99 0 1 6624
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_5
timestamp 1763765945
transform -1 0 99 0 1 9048
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_6
timestamp 1763765945
transform -1 0 99 0 1 1776
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_7
timestamp 1763765945
transform -1 0 99 0 1 4200
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_8
timestamp 1763765945
transform -1 0 99 0 1 564
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_9
timestamp 1763765945
transform -1 0 99 0 1 19956
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_10
timestamp 1763765945
transform -1 0 99 0 1 23592
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_11
timestamp 1763765945
transform -1 0 99 0 1 22380
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_12
timestamp 1763765945
transform -1 0 99 0 1 24804
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_13
timestamp 1763765945
transform -1 0 99 0 1 21168
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_14
timestamp 1763765945
transform -1 0 99 0 1 12684
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_15
timestamp 1763765945
transform -1 0 99 0 1 17532
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_16
timestamp 1763765945
transform -1 0 99 0 1 15108
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_17
timestamp 1763765945
transform -1 0 99 0 1 16320
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_18
timestamp 1763765945
transform -1 0 99 0 1 18744
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_19
timestamp 1763765945
transform -1 0 99 0 1 13896
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_20
timestamp 1763765945
transform -1 0 99 0 1 28440
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_21
timestamp 1763765945
transform -1 0 99 0 1 30864
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_22
timestamp 1763765945
transform -1 0 99 0 1 33288
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_23
timestamp 1763765945
transform -1 0 99 0 1 38136
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_24
timestamp 1763765945
transform -1 0 99 0 1 35712
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_25
timestamp 1763765945
transform -1 0 99 0 1 27228
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_26
timestamp 1763765945
transform -1 0 99 0 1 29652
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_27
timestamp 1763765945
transform -1 0 99 0 1 32076
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_28
timestamp 1763765945
transform -1 0 99 0 1 36924
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_29
timestamp 1763765945
transform -1 0 99 0 1 34500
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_30
timestamp 1763765945
transform -1 0 99 0 1 26016
box 62 103 538 1445
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_31
timestamp 1763765945
transform -1 0 99 0 1 11472
box 62 103 538 1445
use 018SRAM_cell1_512x8m81  018SRAM_cell1_512x8m81_0
timestamp 1763765945
transform -1 0 99 0 1 0
box 62 89 538 797
use 018SRAM_cell1_512x8m81  018SRAM_cell1_512x8m81_1
timestamp 1763765945
transform -1 0 99 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_0
timestamp 1763765945
transform -1 0 11822 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_1
timestamp 1763765945
transform -1 0 11386 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_2
timestamp 1763765945
transform -1 0 10950 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_3
timestamp 1763765945
transform -1 0 10514 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_4
timestamp 1763765945
transform -1 0 9642 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_5
timestamp 1763765945
transform -1 0 10078 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_6
timestamp 1763765945
transform -1 0 9206 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_7
timestamp 1763765945
transform -1 0 8770 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_8
timestamp 1763765945
transform -1 0 12678 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_9
timestamp 1763765945
transform -1 0 13114 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_10
timestamp 1763765945
transform -1 0 13986 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_11
timestamp 1763765945
transform -1 0 13550 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_12
timestamp 1763765945
transform -1 0 14422 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_13
timestamp 1763765945
transform -1 0 14858 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_14
timestamp 1763765945
transform -1 0 15294 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_15
timestamp 1763765945
transform -1 0 15730 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_16
timestamp 1763765945
transform -1 0 5298 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_17
timestamp 1763765945
transform -1 0 6170 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_18
timestamp 1763765945
transform -1 0 5734 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_19
timestamp 1763765945
transform -1 0 6606 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_20
timestamp 1763765945
transform -1 0 7042 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_21
timestamp 1763765945
transform -1 0 7478 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_22
timestamp 1763765945
transform -1 0 7914 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_23
timestamp 1763765945
transform -1 0 4006 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_24
timestamp 1763765945
transform -1 0 3570 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_25
timestamp 1763765945
transform -1 0 3134 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_26
timestamp 1763765945
transform -1 0 2698 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_27
timestamp 1763765945
transform -1 0 1826 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_28
timestamp 1763765945
transform -1 0 2262 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_29
timestamp 1763765945
transform -1 0 1390 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_30
timestamp 1763765945
transform -1 0 954 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_31
timestamp 1763765945
transform -1 0 4862 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_32
timestamp 1763765945
transform -1 0 2698 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_33
timestamp 1763765945
transform -1 0 1826 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_34
timestamp 1763765945
transform -1 0 2262 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_35
timestamp 1763765945
transform -1 0 1390 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_36
timestamp 1763765945
transform -1 0 954 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_37
timestamp 1763765945
transform -1 0 3570 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_38
timestamp 1763765945
transform -1 0 3134 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_39
timestamp 1763765945
transform -1 0 7478 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_40
timestamp 1763765945
transform -1 0 4862 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_41
timestamp 1763765945
transform -1 0 7914 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_42
timestamp 1763765945
transform -1 0 5298 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_43
timestamp 1763765945
transform -1 0 6170 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_44
timestamp 1763765945
transform -1 0 5734 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_45
timestamp 1763765945
transform -1 0 6606 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_46
timestamp 1763765945
transform -1 0 7042 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_47
timestamp 1763765945
transform -1 0 4006 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_48
timestamp 1763765945
transform -1 0 9642 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_49
timestamp 1763765945
transform -1 0 11386 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_50
timestamp 1763765945
transform -1 0 8770 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_51
timestamp 1763765945
transform -1 0 9206 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_52
timestamp 1763765945
transform -1 0 11822 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_53
timestamp 1763765945
transform -1 0 10078 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_54
timestamp 1763765945
transform -1 0 10514 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_55
timestamp 1763765945
transform -1 0 10950 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_56
timestamp 1763765945
transform -1 0 13550 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_57
timestamp 1763765945
transform -1 0 13114 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_59
timestamp 1763765945
transform -1 0 14422 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_60
timestamp 1763765945
transform -1 0 15294 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_61
timestamp 1763765945
transform -1 0 13986 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_62
timestamp 1763765945
transform -1 0 15730 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_63
timestamp 1763765945
transform -1 0 12678 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_64
timestamp 1763765945
transform -1 0 14858 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_0
timestamp 1763765945
transform 1 0 15986 0 -1 5100
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_1
timestamp 1763765945
transform 1 0 15986 0 -1 6312
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_2
timestamp 1763765945
transform 1 0 15986 0 -1 3888
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_3
timestamp 1763765945
transform 1 0 15986 0 -1 2676
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_4
timestamp 1763765945
transform 1 0 15986 0 -1 7524
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_5
timestamp 1763765945
transform 1 0 15986 0 -1 12372
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_6
timestamp 1763765945
transform 1 0 15986 0 -1 11160
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_7
timestamp 1763765945
transform 1 0 15986 0 -1 9948
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_8
timestamp 1763765945
transform 1 0 15986 0 -1 8736
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_9
timestamp 1763765945
transform 1 0 15986 0 -1 1464
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_10
timestamp 1763765945
transform 1 0 15986 0 1 3636
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_11
timestamp 1763765945
transform 1 0 15986 0 1 4848
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_12
timestamp 1763765945
transform 1 0 15986 0 1 7272
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_13
timestamp 1763765945
transform 1 0 15986 0 1 9696
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_14
timestamp 1763765945
transform 1 0 15986 0 1 2424
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_15
timestamp 1763765945
transform 1 0 15986 0 1 6060
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_16
timestamp 1763765945
transform 1 0 15986 0 1 8484
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_17
timestamp 1763765945
transform 1 0 15986 0 1 10908
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_18
timestamp 1763765945
transform 1 0 15986 0 1 1212
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_19
timestamp 1763765945
transform 1 0 15986 0 1 0
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_20
timestamp 1763765945
transform 1 0 15986 0 -1 25704
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_21
timestamp 1763765945
transform 1 0 15986 0 -1 20856
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_22
timestamp 1763765945
transform 1 0 15986 0 -1 24492
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_23
timestamp 1763765945
transform 1 0 15986 0 -1 23280
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_24
timestamp 1763765945
transform 1 0 15986 0 -1 22068
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_25
timestamp 1763765945
transform 1 0 15986 0 -1 16008
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_26
timestamp 1763765945
transform 1 0 15986 0 -1 13584
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_27
timestamp 1763765945
transform 1 0 15986 0 -1 14796
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_28
timestamp 1763765945
transform 1 0 15986 0 -1 19644
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_29
timestamp 1763765945
transform 1 0 15986 0 -1 18432
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_30
timestamp 1763765945
transform 1 0 15986 0 -1 17220
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_31
timestamp 1763765945
transform 1 0 15986 0 1 24240
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_32
timestamp 1763765945
transform 1 0 15986 0 1 20604
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_33
timestamp 1763765945
transform 1 0 15986 0 1 14544
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_34
timestamp 1763765945
transform 1 0 15986 0 1 16968
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_35
timestamp 1763765945
transform 1 0 15986 0 1 19392
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_36
timestamp 1763765945
transform 1 0 15986 0 1 21816
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_37
timestamp 1763765945
transform 1 0 15986 0 1 23028
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_38
timestamp 1763765945
transform 1 0 15986 0 1 13332
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_39
timestamp 1763765945
transform 1 0 15986 0 1 15756
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_40
timestamp 1763765945
transform 1 0 15986 0 1 18180
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_41
timestamp 1763765945
transform 1 0 15986 0 1 25452
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_42
timestamp 1763765945
transform 1 0 15986 0 -1 37824
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_43
timestamp 1763765945
transform 1 0 15986 0 -1 35400
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_44
timestamp 1763765945
transform 1 0 15986 0 -1 32976
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_45
timestamp 1763765945
transform 1 0 15986 0 -1 29340
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_46
timestamp 1763765945
transform 1 0 15986 0 -1 28128
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_47
timestamp 1763765945
transform 1 0 15986 0 -1 39036
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_48
timestamp 1763765945
transform 1 0 15986 0 -1 36612
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_49
timestamp 1763765945
transform 1 0 15986 0 -1 34188
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_50
timestamp 1763765945
transform 1 0 15986 0 -1 31764
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_51
timestamp 1763765945
transform 1 0 15986 0 -1 30552
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_52
timestamp 1763765945
transform 1 0 15986 0 -1 40248
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_53
timestamp 1763765945
transform 1 0 15986 0 1 36360
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_54
timestamp 1763765945
transform 1 0 15986 0 1 26664
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_55
timestamp 1763765945
transform 1 0 15986 0 1 31512
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_56
timestamp 1763765945
transform 1 0 15986 0 1 37572
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_57
timestamp 1763765945
transform 1 0 15986 0 1 33936
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_58
timestamp 1763765945
transform 1 0 15986 0 1 29088
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_59
timestamp 1763765945
transform 1 0 15986 0 1 38784
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_60
timestamp 1763765945
transform 1 0 15986 0 1 30300
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_61
timestamp 1763765945
transform 1 0 15986 0 1 35148
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_62
timestamp 1763765945
transform 1 0 15986 0 1 27876
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_63
timestamp 1763765945
transform 1 0 15986 0 1 32724
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_64
timestamp 1763765945
transform 1 0 15986 0 -1 26916
box 62 89 538 797
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_65
timestamp 1763765945
transform 1 0 15986 0 1 12120
box 62 89 538 797
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_0
timestamp 1763765945
transform -1 0 12251 0 1 0
box 91 55 511 797
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_1
timestamp 1763765945
transform -1 0 4435 0 1 0
box 91 55 511 797
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_2
timestamp 1763765945
transform -1 0 527 0 1 0
box 91 55 511 797
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_3
timestamp 1763765945
transform -1 0 4435 0 -1 40248
box 91 55 511 797
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_4
timestamp 1763765945
transform -1 0 12251 0 -1 40248
box 91 55 511 797
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_5
timestamp 1763765945
transform 1 0 15557 0 -1 40248
box 91 55 511 797
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_6
timestamp 1763765945
transform -1 0 8343 0 1 0
box 91 55 511 797
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_7
timestamp 1763765945
transform -1 0 8343 0 -1 40248
box 91 55 511 797
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_0
timestamp 1763765945
transform 1 0 15557 0 1 0
box 91 55 511 797
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_54
timestamp 1763765945
transform -1 0 527 0 -1 40248
box 91 55 511 797
use M1_NWELL$$44998700_512x8m81  M1_NWELL$$44998700_512x8m81_0
timestamp 1763765945
transform 1 0 16322 0 1 -14699
box -154 -159 154 159
use M1_NWELL$$44998700_512x8m81  M1_NWELL$$44998700_512x8m81_1
timestamp 1763765945
transform 1 0 15941 0 1 -14699
box -154 -159 154 159
use M1_NWELL$$46277676_512x8m81  M1_NWELL$$46277676_512x8m81_0
timestamp 1763765945
transform 1 0 16135 0 1 -9455
box -265 -159 265 159
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_0
timestamp 1763765945
transform 1 0 16620 0 -1 4974
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_1
timestamp 1763765945
transform 1 0 16620 0 -1 3762
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_2
timestamp 1763765945
transform 1 0 16620 0 -1 1338
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_3
timestamp 1763765945
transform 1 0 16620 0 -1 126
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_4
timestamp 1763765945
transform 1 0 16620 0 -1 11034
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_5
timestamp 1763765945
transform 1 0 16620 0 -1 8610
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_6
timestamp 1763765945
transform 1 0 16620 0 -1 6186
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_7
timestamp 1763765945
transform 1 0 16620 0 -1 9822
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_8
timestamp 1763765945
transform 1 0 16620 0 -1 7398
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_9
timestamp 1763765945
transform 1 0 16620 0 -1 2550
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_10
timestamp 1763765945
transform 1 0 16620 0 -1 14670
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_11
timestamp 1763765945
transform 1 0 16620 0 -1 25578
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_12
timestamp 1763765945
transform 1 0 16620 0 -1 24366
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_13
timestamp 1763765945
transform 1 0 16620 0 -1 23154
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_14
timestamp 1763765945
transform 1 0 16620 0 -1 21942
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_15
timestamp 1763765945
transform 1 0 16620 0 -1 20730
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_16
timestamp 1763765945
transform 1 0 16620 0 -1 18306
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_17
timestamp 1763765945
transform 1 0 16620 0 -1 15882
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_18
timestamp 1763765945
transform 1 0 16620 0 -1 13458
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_19
timestamp 1763765945
transform 1 0 16620 0 -1 19518
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_20
timestamp 1763765945
transform 1 0 16620 0 -1 17094
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_21
timestamp 1763765945
transform 1 0 16620 0 -1 37698
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_22
timestamp 1763765945
transform 1 0 16620 0 -1 36486
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_23
timestamp 1763765945
transform 1 0 16620 0 -1 35274
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_24
timestamp 1763765945
transform 1 0 16620 0 -1 34062
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_25
timestamp 1763765945
transform 1 0 16620 0 -1 32850
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_26
timestamp 1763765945
transform 1 0 16620 0 -1 31638
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_27
timestamp 1763765945
transform 1 0 16620 0 -1 30426
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_28
timestamp 1763765945
transform 1 0 16620 0 -1 29214
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_29
timestamp 1763765945
transform 1 0 16620 0 -1 28002
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_30
timestamp 1763765945
transform 1 0 16620 0 -1 26790
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_31
timestamp 1763765945
transform 1 0 16620 0 -1 38910
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_32
timestamp 1763765945
transform 1 0 16620 0 -1 40122
box -96 -124 67 124
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_33
timestamp 1763765945
transform 1 0 16620 0 -1 12246
box -96 -124 67 124
use M1_POLY2$$46559276_512x8m81_0  M1_POLY2$$46559276_512x8m81_0_0
timestamp 1763765945
transform -1 0 15966 0 1 -12400
box -123 -48 123 48
use M1_POLY2$$46559276_512x8m81_0  M1_POLY2$$46559276_512x8m81_0_1
timestamp 1763765945
transform 1 0 16375 0 1 -10338
box -123 -48 123 48
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_0
timestamp 1763765945
transform 1 0 -499 0 1 128
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_1
timestamp 1763765945
transform 1 0 -499 0 1 1340
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_2
timestamp 1763765945
transform 1 0 -499 0 1 2552
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_3
timestamp 1763765945
transform 1 0 -499 0 1 4976
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_4
timestamp 1763765945
transform 1 0 -499 0 1 3764
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_5
timestamp 1763765945
transform 1 0 -499 0 1 9824
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_6
timestamp 1763765945
transform 1 0 -499 0 1 8612
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_7
timestamp 1763765945
transform 1 0 -499 0 1 11036
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_8
timestamp 1763765945
transform 1 0 -499 0 1 12248
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_9
timestamp 1763765945
transform 1 0 -499 0 1 7400
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_10
timestamp 1763765945
transform 1 0 -499 0 1 6188
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_11
timestamp 1763765945
transform 1 0 -499 0 1 14672
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_12
timestamp 1763765945
transform 1 0 -499 0 1 13460
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_13
timestamp 1763765945
transform 1 0 -499 0 1 15884
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_14
timestamp 1763765945
transform 1 0 -499 0 1 17096
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_15
timestamp 1763765945
transform 1 0 -499 0 1 19520
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_16
timestamp 1763765945
transform 1 0 -499 0 1 18308
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_17
timestamp 1763765945
transform 1 0 -499 0 1 20732
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_18
timestamp 1763765945
transform 1 0 -499 0 1 21944
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_19
timestamp 1763765945
transform 1 0 -499 0 1 24368
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_20
timestamp 1763765945
transform 1 0 -499 0 1 23156
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_21
timestamp 1763765945
transform 1 0 -499 0 1 25580
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_22
timestamp 1763765945
transform 1 0 -499 0 1 26792
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_23
timestamp 1763765945
transform 1 0 -499 0 1 29216
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_24
timestamp 1763765945
transform 1 0 -499 0 1 28004
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_25
timestamp 1763765945
transform 1 0 -499 0 1 30428
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_26
timestamp 1763765945
transform 1 0 -499 0 1 31640
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_27
timestamp 1763765945
transform 1 0 -499 0 1 34064
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_28
timestamp 1763765945
transform 1 0 -499 0 1 32852
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_29
timestamp 1763765945
transform 1 0 -499 0 1 35276
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_30
timestamp 1763765945
transform 1 0 -499 0 1 36488
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_31
timestamp 1763765945
transform 1 0 -499 0 1 38912
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_32
timestamp 1763765945
transform 1 0 -499 0 1 37700
box -36 -80 36 78
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_33
timestamp 1763765945
transform 1 0 -499 0 1 40124
box -36 -80 36 78
use M1_PSUB$$46274604_512x8m81  M1_PSUB$$46274604_512x8m81_0
timestamp 1763765945
transform 1 0 16174 0 1 -10851
box -166 -58 166 58
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1763765945
transform 1 0 16618 0 -1 11034
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_1
timestamp 1763765945
transform 1 0 16618 0 -1 8610
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_2
timestamp 1763765945
transform 1 0 16618 0 -1 6185
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_3
timestamp 1763765945
transform 1 0 16618 0 -1 3761
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_4
timestamp 1763765945
transform 1 0 16618 0 -1 1339
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_5
timestamp 1763765945
transform 1 0 16618 0 -1 7398
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_6
timestamp 1763765945
transform 1 0 16618 0 -1 2550
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_7
timestamp 1763765945
transform 1 0 16618 0 -1 127
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_8
timestamp 1763765945
transform 1 0 16618 0 -1 9825
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_9
timestamp 1763765945
transform 1 0 16618 0 -1 4974
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_10
timestamp 1763765945
transform 1 0 16618 0 -1 21942
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_11
timestamp 1763765945
transform 1 0 16618 0 -1 20730
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_12
timestamp 1763765945
transform 1 0 16618 0 -1 18306
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_13
timestamp 1763765945
transform 1 0 16618 0 -1 15882
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_14
timestamp 1763765945
transform 1 0 16618 0 -1 13458
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_15
timestamp 1763765945
transform 1 0 16618 0 -1 17097
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_16
timestamp 1763765945
transform 1 0 16618 0 -1 19518
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_17
timestamp 1763765945
transform 1 0 16618 0 -1 25578
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_18
timestamp 1763765945
transform 1 0 16618 0 -1 14673
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_19
timestamp 1763765945
transform 1 0 16618 0 -1 24366
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_20
timestamp 1763765945
transform 1 0 16618 0 -1 23154
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_21
timestamp 1763765945
transform 1 0 16618 0 -1 37698
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_22
timestamp 1763765945
transform 1 0 16618 0 -1 36486
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_23
timestamp 1763765945
transform 1 0 16618 0 -1 35274
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_24
timestamp 1763765945
transform 1 0 16618 0 -1 34062
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_25
timestamp 1763765945
transform 1 0 16618 0 -1 32850
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_26
timestamp 1763765945
transform 1 0 16618 0 -1 31638
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_27
timestamp 1763765945
transform 1 0 16618 0 -1 30426
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_28
timestamp 1763765945
transform 1 0 16618 0 -1 29214
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_29
timestamp 1763765945
transform 1 0 16618 0 -1 28002
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_30
timestamp 1763765945
transform 1 0 16618 0 -1 26790
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_31
timestamp 1763765945
transform 1 0 16618 0 -1 40122
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_32
timestamp 1763765945
transform 1 0 16618 0 -1 38910
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_33
timestamp 1763765945
transform 1 0 16618 0 -1 12249
box -43 -122 43 122
use M2_M1$$47117356_512x8m81  M2_M1$$47117356_512x8m81_0
timestamp 1763765945
transform 1 0 16179 0 1 -13308
box -45 -1474 45 1874
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_0
timestamp 1763765945
transform 1 0 -499 0 1 1340
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_1
timestamp 1763765945
transform 1 0 -499 0 1 2552
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_2
timestamp 1763765945
transform 1 0 -499 0 1 3764
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_3
timestamp 1763765945
transform 1 0 -499 0 1 4976
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_4
timestamp 1763765945
transform 1 0 -499 0 1 6188
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_5
timestamp 1763765945
transform 1 0 -499 0 1 7400
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_6
timestamp 1763765945
transform 1 0 -499 0 1 8612
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_7
timestamp 1763765945
transform 1 0 -499 0 1 9824
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_8
timestamp 1763765945
transform 1 0 -499 0 1 11036
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_9
timestamp 1763765945
transform 1 0 -499 0 1 12248
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_10
timestamp 1763765945
transform 1 0 -499 0 1 25580
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_11
timestamp 1763765945
transform 1 0 -499 0 1 24368
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_12
timestamp 1763765945
transform 1 0 -499 0 1 23156
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_13
timestamp 1763765945
transform 1 0 -499 0 1 21944
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_14
timestamp 1763765945
transform 1 0 -499 0 1 20732
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_15
timestamp 1763765945
transform 1 0 -499 0 1 19520
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_16
timestamp 1763765945
transform 1 0 -499 0 1 18308
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_17
timestamp 1763765945
transform 1 0 -499 0 1 17096
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_18
timestamp 1763765945
transform 1 0 -499 0 1 13460
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_19
timestamp 1763765945
transform 1 0 -499 0 1 14672
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_20
timestamp 1763765945
transform 1 0 -502 0 1 15884
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_21
timestamp 1763765945
transform 1 0 -499 0 1 38911
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_22
timestamp 1763765945
transform 1 0 -499 0 1 37700
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_23
timestamp 1763765945
transform 1 0 -499 0 1 36488
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_24
timestamp 1763765945
transform 1 0 -499 0 1 35276
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_25
timestamp 1763765945
transform 1 0 -499 0 1 34063
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_26
timestamp 1763765945
transform 1 0 -499 0 1 32852
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_27
timestamp 1763765945
transform 1 0 -499 0 1 31640
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_28
timestamp 1763765945
transform 1 0 -499 0 1 30428
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_29
timestamp 1763765945
transform 1 0 -499 0 1 29216
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_30
timestamp 1763765945
transform 1 0 -499 0 1 28004
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_31
timestamp 1763765945
transform 1 0 -499 0 1 26792
box -34 -99 34 99
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_32
timestamp 1763765945
transform 1 0 -499 0 1 40081
box -34 -99 34 99
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_0
timestamp 1763765945
transform 0 -1 -532 1 0 128
box -35 -99 35 99
use nmos_5p04310591302096_512x8m81  nmos_5p04310591302096_512x8m81_0
timestamp 1763765945
transform 1 0 16098 0 1 -12302
box -116 -44 276 837
use nmos_5p04310591302098_512x8m81  nmos_5p04310591302098_512x8m81_0
timestamp 1763765945
transform 1 0 16095 0 1 -10642
box -116 -44 276 172
use pmos_5p04310591302095_512x8m81  pmos_5p04310591302095_512x8m81_0
timestamp 1763765945
transform 1 0 16095 0 1 -10236
box -202 -86 362 413
use pmos_5p04310591302097_512x8m81  pmos_5p04310591302097_512x8m81_0
timestamp 1763765945
transform 1 0 16098 0 -1 -12498
box -202 -86 362 1079
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_0
timestamp 1763765945
transform 1 0 16298 0 1 -11832
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_1
timestamp 1763765945
transform 1 0 16299 0 1 -10049
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_2
timestamp 1763765945
transform 1 0 16301 0 1 -14577
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_3
timestamp 1763765945
transform 1 0 15992 0 1 -14297
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_4
timestamp 1763765945
transform 1 0 15989 0 1 -11456
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_5
timestamp 1763765945
transform 1 0 15989 0 1 -12256
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_6
timestamp 1763765945
transform 1 0 15985 0 1 -10049
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_7
timestamp 1763765945
transform 1 0 16301 0 1 -14297
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_8
timestamp 1763765945
transform 1 0 15989 0 1 -11832
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_9
timestamp 1763765945
transform 1 0 15992 0 1 -14577
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_10
timestamp 1763765945
transform 1 0 16298 0 1 -11456
box -9 0 73 215
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_11
timestamp 1763765945
transform 1 0 16298 0 1 -12256
box -9 0 73 215
use via1_2_x2_R90_512x8m81_0  via1_2_x2_R90_512x8m81_0_0
timestamp 1763765945
transform 0 -1 16230 1 0 -9489
box -9 0 73 215
use via1_2_x2_R270_512x8m81_0  via1_2_x2_R270_512x8m81_0_0
timestamp 1763765945
transform 0 1 15995 -1 0 -7358
box -9 0 75 215
use ypass_gate_512x8m81_0  ypass_gate_512x8m81_0_0
timestamp 1763765945
transform -1 0 16476 0 1 -9333
box -155 914 651 8659
<< end >>
