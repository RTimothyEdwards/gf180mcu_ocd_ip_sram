magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< psubdiff >>
rect -54 23 1271 56
rect -54 -23 -23 23
rect 1240 -23 1271 23
rect -54 -56 1271 -23
<< psubdiffcont >>
rect -23 -23 1240 23
<< metal1 >>
rect -40 23 1257 42
rect -40 -23 -23 23
rect 1240 -23 1257 23
rect -40 -42 1257 -23
<< end >>
