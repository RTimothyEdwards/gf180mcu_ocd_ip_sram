magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< psubdiff >>
rect -54 23 275 56
rect -54 -23 -23 23
rect 244 -23 275 23
rect -54 -56 275 -23
<< psubdiffcont >>
rect -23 -23 244 23
<< metal1 >>
rect -40 23 261 42
rect -40 -23 -23 23
rect 244 -23 261 23
rect -40 -42 261 -23
<< end >>
