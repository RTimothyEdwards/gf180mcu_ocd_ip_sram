magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal2 >>
rect -266 248 266 275
rect -266 -248 -241 248
rect 241 -248 266 248
rect -266 -275 266 -248
<< via2 >>
rect -241 -248 241 248
<< metal3 >>
rect -266 248 266 275
rect -266 -248 -241 248
rect 241 -248 266 248
rect -266 -275 266 -248
<< end >>
