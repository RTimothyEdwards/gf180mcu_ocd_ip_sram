magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< nwell >>
rect -174 -86 230 1906
<< pmos >>
rect 0 0 56 1820
<< pdiff >>
rect -88 1807 0 1820
rect -88 13 -75 1807
rect -29 13 0 1807
rect -88 0 0 13
rect 56 1807 144 1820
rect 56 13 85 1807
rect 131 13 144 1807
rect 56 0 144 13
<< pdiffc >>
rect -75 13 -29 1807
rect 85 13 131 1807
<< polysilicon >>
rect 0 1820 56 1864
rect 0 -44 56 0
<< metal1 >>
rect -75 1807 -29 1820
rect -75 0 -29 13
rect 85 1807 131 1820
rect 85 0 131 13
<< labels >>
flabel pdiffc -40 910 -40 910 0 FreeSans 186 0 0 0 S
flabel pdiffc 96 910 96 910 0 FreeSans 186 0 0 0 D
<< end >>
