magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< nwell >>
rect 82 512 518 797
<< pwell >>
rect 82 89 518 512
<< sramnfet >>
rect 192 342 248 432
rect 352 342 408 432
rect 110 178 166 250
rect 434 178 490 250
<< srampfet >>
rect 192 592 248 648
rect 352 592 408 648
<< sramndiff >>
rect 110 413 192 432
rect 110 367 117 413
rect 163 367 192 413
rect 110 342 192 367
rect 248 342 352 432
rect 408 413 490 432
rect 408 367 437 413
rect 483 367 490 413
rect 408 342 490 367
rect 110 250 166 342
rect 270 327 330 342
rect 270 281 277 327
rect 323 281 330 327
rect 270 270 330 281
rect 434 250 490 342
rect 110 156 166 178
rect 434 156 490 178
rect 110 149 170 156
rect 110 103 117 149
rect 163 103 170 149
rect 110 96 170 103
rect 430 149 490 156
rect 430 103 437 149
rect 483 103 490 149
rect 430 96 490 103
<< srampdiff >>
rect 270 755 330 766
rect 270 709 277 755
rect 323 709 330 755
rect 110 648 170 654
rect 270 648 330 709
rect 430 648 490 654
rect 110 647 192 648
rect 110 601 117 647
rect 163 601 192 647
rect 110 592 192 601
rect 248 592 352 648
rect 408 647 490 648
rect 408 601 437 647
rect 483 601 490 647
rect 408 592 490 601
<< sramndc >>
rect 117 367 163 413
rect 437 367 483 413
rect 277 281 323 327
rect 117 103 163 149
rect 437 103 483 149
<< srampdc >>
rect 277 709 323 755
rect 117 601 163 647
rect 437 601 483 647
<< polysilicon >>
rect 192 648 248 692
rect 352 648 408 692
rect 192 524 248 592
rect 352 572 408 592
rect 330 559 408 572
rect 192 511 271 524
rect 192 465 212 511
rect 258 465 271 511
rect 330 513 343 559
rect 389 513 408 559
rect 330 500 408 513
rect 192 452 271 465
rect 192 432 248 452
rect 352 432 408 500
rect 192 298 248 342
rect 352 298 408 342
rect 62 178 110 250
rect 166 178 434 250
rect 490 178 538 250
<< polycontact >>
rect 212 465 258 511
rect 343 513 389 559
<< metal1 >>
rect 82 755 518 771
rect 82 709 277 755
rect 323 709 518 755
rect 82 693 518 709
rect 163 601 389 647
rect 117 597 389 601
rect 117 413 166 597
rect 332 559 389 597
rect 163 367 166 413
rect 212 511 268 530
rect 258 465 268 511
rect 332 513 343 559
rect 332 494 389 513
rect 435 601 437 647
rect 212 448 268 465
rect 435 448 483 601
rect 212 413 483 448
rect 212 402 437 413
rect 435 367 437 402
rect 252 327 348 356
rect 252 321 277 327
rect 82 281 277 321
rect 323 321 348 327
rect 323 281 518 321
rect 82 199 518 281
rect 112 149 258 152
rect 112 103 117 149
rect 163 103 258 149
rect 112 100 258 103
rect 342 149 488 152
rect 342 103 437 149
rect 483 103 488 149
rect 342 100 488 103
<< metal2 >>
rect 134 89 254 771
rect 346 89 466 771
<< metal3 >>
rect 82 330 518 690
<< properties >>
string FIXED_BBOX 82 126 518 732
string MASKHINTS_SRAMDEF 82 89 518 797
<< end >>
