magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< psubdiff >>
rect -110 23 111 57
rect -110 -23 -78 23
rect 78 -23 111 23
rect -110 -58 111 -23
<< psubdiffcont >>
rect -78 -23 78 23
<< metal1 >>
rect -105 23 105 51
rect -105 -23 -78 23
rect 78 -23 105 23
rect -105 -51 105 -23
<< end >>
