magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< polysilicon >>
rect -125 -34 -70 0
rect 34 -34 89 0
rect 195 -34 251 0
rect 355 -34 410 0
rect 516 -34 572 0
use nmos_5p04310591302085_3v1024x8m81  nmos_5p04310591302085_3v1024x8m81_0
timestamp 1764525316
transform 1 0 -14 0 1 0
box -200 -44 674 975
<< end >>
