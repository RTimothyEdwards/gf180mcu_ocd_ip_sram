magic
tech gf180mcuD
magscale 1 10
timestamp 1765475971
<< ndiff >>
rect -53 60 53 93
rect -53 -60 -23 60
rect 23 -60 53 60
rect -53 -92 53 -60
<< ndiffc >>
rect -23 -60 23 60
<< metal1 >>
rect -40 60 40 79
rect -40 34 -23 60
rect -53 31 -23 34
rect 23 34 40 60
rect 23 31 53 34
rect -53 -31 -31 31
rect 30 -31 53 31
rect -53 -34 -23 -31
rect -40 -60 -23 -34
rect 23 -34 53 -31
rect 23 -60 40 -34
rect -40 -79 40 -60
<< via1 >>
rect -31 -31 -23 31
rect -23 -31 23 31
rect 23 -31 30 31
<< metal2 >>
rect -43 31 42 34
rect -43 -31 -31 31
rect 30 -31 42 31
rect -43 -34 42 -31
<< end >>
