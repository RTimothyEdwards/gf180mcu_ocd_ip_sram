magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect -928 -501 928 501
<< nsubdiff >>
rect -829 359 829 399
rect -829 -359 -791 359
rect 791 -359 829 359
rect -829 -399 829 -359
<< nsubdiffcont >>
rect -791 -359 791 359
<< metal1 >>
rect -815 359 815 385
rect -815 -359 -791 359
rect 791 -359 815 359
rect -815 -385 815 -359
<< end >>
