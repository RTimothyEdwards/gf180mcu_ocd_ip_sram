magic
tech gf180mcuD
magscale 1 10
timestamp 1764700137
<< metal2 >>
rect 0 196 65 222
rect 0 26 3 196
rect 60 26 65 196
rect 0 0 65 26
<< via2 >>
rect 3 26 60 196
<< metal3 >>
rect -9 196 74 222
rect -9 26 3 196
rect 60 26 74 196
rect -9 0 74 26
<< end >>
