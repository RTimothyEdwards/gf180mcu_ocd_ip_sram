magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< polysilicon >>
rect -14 317 41 351
rect -14 -34 41 0
use nmos_5p04310591302015_512x8m81  nmos_5p04310591302015_512x8m81_0
timestamp 1763765945
transform 1 0 -14 0 1 0
box -88 -44 144 362
<< end >>
