magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nwell >>
rect -320 -159 320 159
<< nsubdiff >>
rect -233 23 244 56
rect -233 -23 -189 23
rect 189 -23 244 23
rect -233 -56 244 -23
<< nsubdiffcont >>
rect -189 -23 189 23
<< metal1 >>
rect -206 23 230 42
rect -206 -23 -189 23
rect 189 -23 230 23
rect -206 -42 230 -23
<< end >>
