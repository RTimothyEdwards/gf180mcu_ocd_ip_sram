magic
tech gf180mcuD
magscale 1 10
timestamp 1763486358
<< nwell >>
rect 441 20127 4028 20391
rect 441 18837 3465 20127
rect 441 17060 4028 18837
rect 3849 17042 4028 17060
rect 225 12681 440 13973
rect 1014 6566 1055 6595
rect 1574 6566 1612 6583
<< metal1 >>
rect 309 18913 373 18974
rect 308 11455 349 11522
rect 3740 7393 3806 8076
rect 1894 6457 1953 6673
rect 2391 5707 2534 5804
rect 1677 979 1729 1053
rect 1842 979 1918 1053
rect 2342 979 2426 1063
rect 1834 603 1918 736
rect 2342 603 2426 736
<< metal2 >>
rect 281 18965 333 18991
rect 277 11488 334 18965
rect 431 11917 487 13545
rect 1280 11991 1336 13449
rect 2197 11991 2259 13464
rect 3101 11992 3164 13460
rect 3878 11844 3934 13520
rect 3544 11780 3934 11844
rect 699 7475 1350 7532
rect 1450 7524 1516 11525
rect 327 345 392 6243
rect 581 5818 648 6565
rect 581 5754 809 5818
rect 742 4465 809 5754
rect 1294 5735 1350 7475
rect 1294 5678 1419 5735
rect 591 4396 809 4465
rect 591 1365 658 4396
rect 1055 4379 1121 4801
rect 1363 4584 1419 5678
rect 1579 5693 1645 11501
rect 1708 7524 1774 11525
rect 2963 6187 3028 6307
rect 3284 6266 3350 6392
rect 3284 6199 3535 6266
rect 2963 6119 3104 6187
rect 3469 6100 3535 6199
rect 1579 5636 1991 5693
rect 935 4292 1121 4379
rect 1310 4527 1419 4584
rect 935 3785 1001 4292
rect 915 3710 1001 3785
rect 591 1240 690 1365
rect 634 230 690 1240
rect 915 1250 981 3710
rect 1310 1651 1366 4527
rect 1589 3837 1647 4446
rect 1924 3877 1991 5636
rect 3740 5067 3806 7478
rect 3740 4997 3826 5067
rect 3076 4481 3300 4575
rect 3760 4541 3826 4997
rect 3239 4262 3300 4481
rect 3587 4473 3826 4541
rect 3587 4262 3645 4473
rect 1495 3798 1647 3837
rect 1736 3821 1991 3877
rect 1736 3598 1802 3821
rect 1579 3513 1802 3598
rect 1579 2671 1645 3513
rect 1310 1598 1380 1651
rect 915 1160 1011 1250
rect 945 340 1011 1160
rect 1319 1034 1380 1598
rect 1319 976 1430 1034
rect 1367 210 1430 976
rect 1367 149 1452 210
rect 1389 -969 1452 149
rect 1389 -1032 2159 -969
rect 2096 -1354 2159 -1032
<< metal3 >>
rect 0 15638 351 17021
rect 263 11544 3861 11704
rect 3845 9438 4055 11344
rect 222 3786 1617 3848
rect 3938 2534 4055 3487
rect 3945 449 4055 767
use din_512x8m81  din_512x8m81_0
timestamp 1763476864
transform 1 0 226 0 1 5808
box -156 -50 1824 6415
use M1_NACTIVE4310591302024_512x8m81  M1_NACTIVE4310591302024_512x8m81_0
timestamp 1763476864
transform 1 0 3909 0 1 600
box -38 -128 36 128
use M2_M1$$45012012_512x8m81  M2_M1$$45012012_512x8m81_0
timestamp 1763476864
transform 1 0 1767 0 1 11654
box -562 -46 562 46
use M2_M1$$45013036_512x8m81  M2_M1$$45013036_512x8m81_0
timestamp 1763476864
transform 1 0 2839 0 1 11654
box -266 -46 266 46
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_0
timestamp 1763476864
transform 0 -1 3614 1 0 4203
box -63 -34 63 34
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_1
timestamp 1763476864
transform 0 -1 3273 1 0 4203
box -63 -34 63 34
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_0
timestamp 1763476864
transform 0 -1 642 1 0 256
box -34 -63 34 63
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_1
timestamp 1763476864
transform 1 0 2126 0 1 -1295
box -34 -63 34 63
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_0
timestamp 1763476864
transform 1 0 299 0 1 18941
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_1
timestamp 1763476864
transform 1 0 461 0 1 13504
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_2
timestamp 1763476864
transform 1 0 3901 0 1 13474
box -35 -56 35 55
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_3
timestamp 1763476864
transform 1 0 307 0 1 11488
box -35 -56 35 55
use M2_M14310591302025_512x8m81  M2_M14310591302025_512x8m81_0
timestamp 1763476864
transform 1 0 3909 0 1 601
box -34 -85 34 135
use m2_saout01_512x8m81  m2_saout01_512x8m81_0
timestamp 1763476864
transform 1 0 480 0 1 20290
box -102 -44 3491 1507
use M3_M2$$43370540_512x8m81  M3_M2$$43370540_512x8m81_0
timestamp 1763476864
transform 1 0 2839 0 1 11654
box -266 -46 266 46
use M3_M2$$44741676_512x8m81  M3_M2$$44741676_512x8m81_0
timestamp 1763476864
transform 1 0 1767 0 1 11654
box -562 -46 562 46
use M3_M2431059130207_512x8m81  M3_M2431059130207_512x8m81_0
timestamp 1763476864
transform 1 0 1554 0 1 3817
box -63 -35 63 35
use M3_M24310591302026_512x8m81  M3_M24310591302026_512x8m81_0
timestamp 1763476864
transform 1 0 3909 0 1 601
box -35 -135 35 135
use mux821_512x8m81  mux821_512x8m81_0
timestamp 1763486358
transform 1 0 387 0 1 12008
box -575 93 4956 8484
use outbuf_oe_512x8m81  outbuf_oe_512x8m81_0
timestamp 1763476864
transform 1 0 442 0 1 4201
box -372 -251 3623 2326
use sa_512x8m81  sa_512x8m81_0
timestamp 1763476864
transform 1 0 442 0 1 6370
box -249 -137 3523 5747
use sacntl_2_512x8m81  sacntl_2_512x8m81_0
timestamp 1763476864
transform 1 0 442 0 1 361
box -371 -16 3623 3958
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_0
timestamp 1763476864
transform 1 0 1451 0 1 8985
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_1
timestamp 1763476864
transform 1 0 1451 0 1 8442
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_2
timestamp 1763476864
transform 1 0 1451 0 1 7801
box -9 0 73 215
use via1_x2_512x8m81  via1_x2_512x8m81_0
timestamp 1763476864
transform -1 0 1644 0 -1 11523
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_1
timestamp 1763476864
transform -1 0 1122 0 -1 4796
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_2
timestamp 1763476864
transform 1 0 1579 0 1 2672
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_3
timestamp 1763476864
transform 1 0 3741 0 1 7317
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_4
timestamp 1763476864
transform 1 0 322 0 1 6116
box -8 0 72 222
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 3592 1 0 11780
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_1
timestamp 1763476864
transform 0 -1 1381 1 0 13456
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_2
timestamp 1763476864
transform 0 -1 2271 1 0 13456
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_3
timestamp 1763476864
transform 0 -1 3185 1 0 13456
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_4
timestamp 1763476864
transform 0 -1 647 1 0 6498
box -8 0 72 215
use via2_512x8m81  via2_512x8m81_0
timestamp 1763476864
transform 1 0 3743 0 1 13431
box 0 0 65 92
use via2_512x8m81  via2_512x8m81_1
timestamp 1763476864
transform 1 0 3135 0 1 13672
box 0 0 65 92
use via2_512x8m81  via2_512x8m81_2
timestamp 1763476864
transform 1 0 2947 0 1 13910
box 0 0 65 92
use via2_512x8m81  via2_512x8m81_3
timestamp 1763476864
transform 1 0 2044 0 1 14695
box 0 0 65 92
use via2_512x8m81  via2_512x8m81_4
timestamp 1763476864
transform 1 0 2229 0 1 14159
box 0 0 65 92
use via2_512x8m81  via2_512x8m81_5
timestamp 1763476864
transform 1 0 1331 0 1 14940
box 0 0 65 92
use via2_512x8m81  via2_512x8m81_6
timestamp 1763476864
transform 1 0 1143 0 1 15181
box 0 0 65 92
use via2_512x8m81  via2_512x8m81_7
timestamp 1763476864
transform 1 0 425 0 1 15404
box 0 0 65 92
use via2_x2_512x8m81  via2_x2_512x8m81_0
timestamp 1763476864
transform 1 0 1709 0 1 8985
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_1
timestamp 1763476864
transform 1 0 1709 0 1 8442
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_2
timestamp 1763476864
transform 1 0 1709 0 1 7801
box -9 0 74 222
use wen_wm1_512x8m81  wen_wm1_512x8m81_0
timestamp 1763486358
transform 1 0 225 0 1 -2018
box -133 -24 3461 2300
<< labels >>
rlabel metal3 s 653 20231 653 20231 4 vdd
port 10 nsew
rlabel metal2 s 3403 20112 3403 20112 4 bb[1]
port 16 nsew
rlabel metal2 s 2682 20115 2682 20115 4 bb[2]
port 18 nsew
rlabel metal2 s 2542 20118 2542 20118 4 bb[3]
port 19 nsew
rlabel metal2 s 1815 20113 1815 20113 4 bb[4]
port 20 nsew
rlabel metal2 s 1670 20113 1670 20113 4 bb[5]
port 21 nsew
rlabel metal2 s 808 20118 808 20118 4 bb[7]
port 22 nsew
rlabel metal2 s 948 20113 948 20113 4 bb[6]
port 23 nsew
rlabel metal2 s 3114 20112 3114 20112 4 b[1]
port 25 nsew
rlabel metal2 s 2104 20112 2104 20112 4 b[4]
port 26 nsew
rlabel metal2 s 1380 20112 1380 20112 4 b[5]
port 27 nsew
rlabel metal2 s 1239 20112 1239 20112 4 b[6]
port 28 nsew
rlabel metal2 s 515 20112 515 20112 4 b[7]
port 29 nsew
rlabel metal2 s 2975 20112 2975 20112 4 b[2]
port 30 nsew
rlabel metal2 s 2247 20112 2247 20112 4 b[3]
port 31 nsew
rlabel metal2 s 511 20112 511 20112 4 b[7]
port 29 nsew
rlabel metal2 s 1237 20112 1237 20112 4 b[6]
port 28 nsew
rlabel metal2 s 1383 20112 1383 20112 4 b[5]
port 27 nsew
rlabel metal2 s 2102 20112 2102 20112 4 b[4]
port 26 nsew
rlabel metal2 s 2245 20112 2245 20112 4 b[3]
port 31 nsew
rlabel metal2 s 2974 20112 2974 20112 4 b[2]
port 30 nsew
rlabel metal2 s 3115 20112 3115 20112 4 b[1]
port 25 nsew
rlabel metal2 s 947 20113 947 20113 4 bb[6]
port 23 nsew
rlabel metal2 s 805 20118 805 20118 4 bb[7]
port 22 nsew
rlabel metal2 s 1673 20113 1673 20113 4 bb[5]
port 21 nsew
rlabel metal2 s 1813 20113 1813 20113 4 bb[4]
port 20 nsew
rlabel metal2 s 2539 20118 2539 20118 4 bb[3]
port 19 nsew
rlabel metal2 s 2679 20115 2679 20115 4 bb[2]
port 18 nsew
rlabel metal2 s 3404 20112 3404 20112 4 bb[1]
port 16 nsew
rlabel metal3 s 616 1366 616 1366 4 men
port 8 nsew
rlabel metal3 s 2042 1103 2042 1103 4 vss
port 9 nsew
rlabel metal3 s 2042 1865 2042 1865 4 vss
port 9 nsew
rlabel metal3 s 567 14482 567 14482 4 ypass[4]
port 4 nsew
rlabel metal3 s 2121 3021 2121 3021 4 vdd
port 10 nsew
rlabel metal3 s 1484 624 1484 624 4 vdd
port 10 nsew
rlabel metal3 s 1957 4169 1957 4169 4 vss
port 9 nsew
rlabel metal3 s 1314 8065 1314 8065 4 vss
port 9 nsew
rlabel metal3 s 567 15153 567 15153 4 ypass[7]
port 7 nsew
rlabel metal3 s 567 14931 567 14931 4 ypass[6]
port 6 nsew
rlabel metal3 s 567 14709 567 14709 4 ypass[5]
port 5 nsew
rlabel metal3 s 567 14023 567 14023 4 ypass[3]
port 3 nsew
rlabel metal3 s 567 13801 567 13801 4 ypass[2]
port 2 nsew
rlabel metal3 s 567 13579 567 13579 4 ypass[1]
port 1 nsew
rlabel metal3 s 664 15750 664 15750 4 vss
port 9 nsew
rlabel metal3 s 653 13054 653 13054 4 vdd
port 10 nsew
rlabel metal3 s 681 12168 681 12168 4 vss
port 9 nsew
rlabel metal3 s 1264 9977 1264 9977 4 vdd
port 10 nsew
rlabel metal3 s 2312 5692 2312 5692 4 vdd
port 10 nsew
rlabel metal3 s 567 13354 567 13354 4 ypass[0]
port 11 nsew
flabel metal3 s 322 -70 322 -70 0 FreeSans 420 0 0 0 VDD
port 12 nsew
flabel metal3 s 322 5308 322 5308 0 FreeSans 420 0 0 0 VDD
port 12 nsew
flabel metal3 s 322 2656 322 2656 0 FreeSans 420 0 0 0 VDD
port 12 nsew
flabel metal3 s 322 655 322 655 0 FreeSans 420 0 0 0 VDD
port 12 nsew
flabel metal3 s 322 -1700 322 -1700 0 FreeSans 420 0 0 0 VDD
port 12 nsew
flabel metal3 s 431 -1059 431 -1059 0 FreeSans 420 0 0 0 GWEN
port 13 nsew
flabel metal3 s 322 2068 322 2068 0 FreeSans 420 0 0 0 VSS
port 14 nsew
flabel metal3 s 322 16697 322 16697 0 FreeSans 420 0 0 0 VSS
port 14 nsew
flabel metal3 s 322 -1231 322 -1231 0 FreeSans 420 0 0 0 VSS
port 14 nsew
flabel metal3 s 322 4768 322 4768 0 FreeSans 420 0 0 0 VSS
port 14 nsew
flabel metal3 s 322 9110 322 9110 0 FreeSans 420 0 0 0 VSS
port 14 nsew
flabel metal3 s 322 -586 322 -586 0 FreeSans 420 0 0 0 VSS
port 14 nsew
flabel metal3 s 322 1096 322 1096 0 FreeSans 420 0 0 0 VSS
port 14 nsew
flabel metal3 s 322 12320 322 12320 0 FreeSans 420 0 0 0 VSS
port 14 nsew
flabel metal3 s 322 -896 322 -896 0 FreeSans 420 0 0 0 VSS
port 14 nsew
flabel metal3 s 322 6315 322 6315 0 FreeSans 420 0 0 0 VDD
port 12 nsew
flabel metal3 s 322 9595 322 9595 0 FreeSans 420 0 0 0 VDD
port 12 nsew
flabel metal3 s 322 12976 322 12976 0 FreeSans 420 0 0 0 VDD
port 12 nsew
flabel metal3 s 450 3816 450 3816 0 FreeSans 420 0 0 0 GWE
port 15 nsew
rlabel metal1 s 695 19297 695 19297 4 pcb
port 34 nsew
rlabel metal1 s 488 6164 488 6164 4 datain
port 32 nsew
rlabel metal1 s 695 19295 695 19295 4 pcb
port 34 nsew
rlabel metal1 s 1260 11499 1260 11499 4 pcb
port 34 nsew
flabel metal1 s 505 -2010 505 -2010 0 FreeSans 420 0 0 0 WEN
port 35 nsew
rlabel metal2 s 975 1131 975 1131 4 q
port 33 nsew
rlabel metal2 s 346 1551 346 1551 4 datain
port 32 nsew
<< end >>
