magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal1 >>
rect -34 127 34 135
rect -34 -77 -26 127
rect 26 -77 34 127
rect -34 -85 34 -77
<< via1 >>
rect -26 -77 26 127
<< metal2 >>
rect -34 127 34 135
rect -34 -77 -26 127
rect 26 -77 34 127
rect -34 -85 34 -77
<< end >>
