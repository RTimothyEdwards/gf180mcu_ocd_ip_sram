magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< error_s >>
rect -117 0 -71 89
rect 43 0 89 89
rect 203 0 249 89
<< nwell >>
rect -133 -65 265 154
<< polysilicon >>
rect -42 89 13 123
rect 118 89 174 123
rect -42 -34 13 0
rect 118 -34 174 0
use pmos_5p0431059130206_3v1024x8m81  pmos_5p0431059130206_3v1024x8m81_0
timestamp 1764525316
transform 1 0 -14 0 1 0
box -202 -86 362 175
<< end >>
