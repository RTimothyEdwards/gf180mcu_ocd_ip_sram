magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
use 018SRAM_strap1_3v512x8m81  018SRAM_strap1_3v512x8m81_0
timestamp 1763765945
transform 1 0 0 0 -1 0
box 91 55 511 797
use 018SRAM_strap1_3v512x8m81  018SRAM_strap1_3v512x8m81_1
timestamp 1763765945
transform 1 0 0 0 1 -252
box 91 55 511 797
<< end >>
