magic
tech gf180mcuD
magscale 1 10
timestamp 1765924077
<< nwell >>
rect -32 10266 602 11861
rect -7 9396 602 10266
rect -5 8409 602 9396
rect -5 4935 633 5208
rect -130 4479 633 4935
<< pmos >>
rect 172 10921 228 11239
rect 332 10921 388 11239
rect 172 10416 228 10733
rect 332 10416 388 10733
rect 169 4568 225 4707
rect 376 4568 432 4707
<< ndiff >>
rect 54 4319 80 4391
rect 489 4319 505 4391
<< pdiff >>
rect 54 11195 172 11239
rect 54 11149 97 11195
rect 143 11149 172 11195
rect 54 11013 172 11149
rect 54 10967 97 11013
rect 143 10967 172 11013
rect 54 10921 172 10967
rect 228 11195 332 11239
rect 228 11149 257 11195
rect 303 11149 332 11195
rect 228 11013 332 11149
rect 228 10967 257 11013
rect 303 10967 332 11013
rect 228 10921 332 10967
rect 388 11195 505 11239
rect 388 11149 419 11195
rect 465 11149 505 11195
rect 388 11013 505 11149
rect 388 10967 419 11013
rect 465 10967 505 11013
rect 388 10921 505 10967
rect 54 10690 172 10733
rect 54 10644 97 10690
rect 143 10644 172 10690
rect 54 10508 172 10644
rect 54 10462 97 10508
rect 143 10462 172 10508
rect 54 10416 172 10462
rect 228 10690 332 10733
rect 228 10644 257 10690
rect 303 10644 332 10690
rect 228 10508 332 10644
rect 228 10462 257 10508
rect 303 10462 332 10508
rect 228 10416 332 10462
rect 388 10690 505 10733
rect 388 10644 419 10690
rect 465 10644 505 10690
rect 388 10508 505 10644
rect 388 10462 419 10508
rect 465 10462 505 10508
rect 388 10416 505 10462
rect 36 4662 169 4707
rect 36 4615 78 4662
rect 124 4615 169 4662
rect 36 4568 169 4615
rect 225 4661 376 4707
rect 225 4615 280 4661
rect 326 4615 376 4661
rect 225 4568 376 4615
rect 432 4661 547 4707
rect 432 4615 482 4661
rect 528 4615 547 4661
rect 432 4568 547 4615
<< pdiffc >>
rect 97 11149 143 11195
rect 97 10967 143 11013
rect 257 11149 303 11195
rect 257 10967 303 11013
rect 419 11149 465 11195
rect 419 10967 465 11013
rect 97 10644 143 10690
rect 97 10462 143 10508
rect 257 10644 303 10690
rect 257 10462 303 10508
rect 419 10644 465 10690
rect 419 10462 465 10508
rect 78 4615 124 4662
rect 280 4615 326 4661
rect 482 4615 528 4661
<< nsubdiff >>
rect 119 11552 516 11712
<< polysilicon >>
rect 172 11239 228 11436
rect 332 11239 388 11436
rect 172 10733 228 10921
rect 332 10733 388 10921
rect 172 10352 228 10416
rect 332 10352 388 10416
rect 172 10268 388 10352
rect 172 10267 304 10268
rect 248 10118 304 10267
rect 250 8479 306 8553
rect 250 8400 315 8479
rect 250 6868 306 7515
rect 250 6045 306 6148
rect 250 5900 306 5952
rect 250 5853 306 5888
rect 169 4846 432 4945
rect 169 4707 225 4846
rect 376 4707 432 4846
rect 169 4518 225 4568
rect 376 4519 432 4568
rect 169 4470 228 4518
rect 172 4425 228 4470
rect 340 4470 432 4519
rect 340 4425 396 4470
rect 172 4257 228 4286
rect 340 4257 396 4286
<< metal1 >>
rect 50 11562 510 11717
rect 77 11434 480 11562
rect 77 11195 159 11434
rect 77 11149 97 11195
rect 143 11149 159 11195
rect 77 11013 159 11149
rect 77 10967 97 11013
rect 143 10967 159 11013
rect 77 10690 159 10967
rect 222 11195 337 11382
rect 222 11149 257 11195
rect 303 11149 337 11195
rect 222 11013 337 11149
rect 222 10967 257 11013
rect 303 10967 337 11013
rect 222 10930 337 10967
rect 402 11195 480 11434
rect 402 11149 419 11195
rect 465 11149 480 11195
rect 402 11013 480 11149
rect 402 10967 419 11013
rect 465 10967 480 11013
rect 77 10644 97 10690
rect 143 10644 159 10690
rect 77 10508 159 10644
rect 77 10462 97 10508
rect 143 10462 159 10508
rect 77 10425 159 10462
rect 222 10690 337 10879
rect 222 10644 257 10690
rect 303 10644 337 10690
rect 222 10508 337 10644
rect 222 10462 257 10508
rect 303 10462 337 10508
rect 222 10425 337 10462
rect 402 10690 480 10967
rect 402 10644 419 10690
rect 465 10644 480 10690
rect 402 10508 480 10644
rect 402 10462 419 10508
rect 465 10462 480 10508
rect 402 10425 480 10462
rect 88 9710 219 9890
rect 333 9710 463 9890
rect 88 9066 182 9240
rect 138 8750 182 9066
rect 119 8673 182 8750
rect 381 9075 463 9240
rect 119 7560 189 8673
rect 239 8296 315 8480
rect 381 7496 465 9075
rect 45 7381 465 7496
rect 43 7103 506 7237
rect 123 6938 329 7035
rect 123 6191 188 6938
rect 380 6233 433 6816
rect 123 5765 180 6191
rect 232 6021 328 6124
rect 227 5873 328 5968
rect 123 5181 181 5765
rect 378 5187 433 6233
rect 54 4662 131 5086
rect 199 4856 329 4953
rect 54 4615 78 4662
rect 124 4615 131 4662
rect 54 4577 131 4615
rect 245 4661 328 4777
rect 245 4615 280 4661
rect 326 4615 328 4661
rect 53 4218 157 4389
rect 245 4327 328 4615
rect 466 4661 537 5086
rect 466 4615 482 4661
rect 528 4615 537 4661
rect 466 4577 537 4615
rect 415 4218 505 4387
rect 53 4096 505 4218
<< metal2 >>
rect 88 11314 144 11715
rect 216 11435 344 11717
rect 245 11434 344 11435
rect 88 11258 327 11314
rect 88 9109 144 11258
rect 421 10808 477 11715
rect 285 10752 477 10808
rect 26 7494 82 7495
rect 26 7424 129 7494
rect 26 4011 82 7424
rect 248 7368 304 8406
rect 138 7312 304 7368
rect 138 5965 194 7312
rect 421 7071 477 10752
rect 250 7015 477 7071
rect 381 6124 444 6953
rect 260 6027 444 6124
rect 138 5938 245 5965
rect 138 5882 312 5938
rect 138 5854 245 5882
rect 138 4777 194 5854
rect 381 5494 444 6027
rect 250 5397 444 5494
rect 250 4846 306 5397
rect 138 4598 326 4777
rect 138 4597 290 4598
rect 172 4063 272 4225
<< metal3 >>
rect -65 10338 525 11716
rect -41 7127 525 8527
rect -41 6881 525 7021
rect -41 6639 525 6779
rect -41 6398 525 6538
rect -41 6156 525 6296
rect -41 5924 525 6064
rect -41 5682 525 5822
rect -41 5440 525 5580
rect -41 5198 525 5338
rect -41 4610 525 5052
rect -41 4017 525 4464
use M1_NWELL05_3v512x8m81  M1_NWELL05_3v512x8m81_0
timestamp 1764525316
transform 1 0 285 0 1 11632
box -265 -159 265 159
use M1_NWELL09_3v512x8m81  M1_NWELL09_3v512x8m81_1
timestamp 1764525316
transform 1 0 287 0 1 5043
box -320 -159 330 159
use M1_POLY24310591302030_3v512x8m81  M1_POLY24310591302030_3v512x8m81_0
timestamp 1764525316
transform 1 0 272 0 1 10310
box -95 -36 95 36
use M1_POLY24310591302031_3v512x8m81  M1_POLY24310591302031_3v512x8m81_0
timestamp 1764525316
transform 1 0 253 0 1 4903
box -36 -36 36 36
use M1_POLY24310591302031_3v512x8m81  M1_POLY24310591302031_3v512x8m81_1
timestamp 1764525316
transform 1 0 280 0 1 5910
box -36 -36 36 36
use M1_POLY24310591302031_3v512x8m81  M1_POLY24310591302031_3v512x8m81_2
timestamp 1764525316
transform 1 0 281 0 1 6087
box -36 -36 36 36
use M1_POLY24310591302031_3v512x8m81  M1_POLY24310591302031_3v512x8m81_6
timestamp 1764525316
transform 1 0 276 0 1 8442
box -36 -36 36 36
use M1_PSUB$$45111340_3v512x8m81  M1_PSUB$$45111340_3v512x8m81_0
timestamp 1764525316
transform 1 0 150 0 1 7168
box -56 -58 56 58
use M1_PSUB$$47122476_3v512x8m81  M1_PSUB$$47122476_3v512x8m81_0
timestamp 1764525316
transform 1 0 277 0 1 4160
box -223 -58 254 57
use M2_M1431059130208_3v512x8m81  M2_M1431059130208_3v512x8m81_0
timestamp 1764525316
transform 1 0 287 0 1 4687
box -34 -63 34 63
use M2_M1431059130208_3v512x8m81  M2_M1431059130208_3v512x8m81_2
timestamp 1764525316
transform 1 0 122 0 1 9800
box -34 -63 34 63
use M2_M1431059130208_3v512x8m81  M2_M1431059130208_3v512x8m81_3
timestamp 1764525316
transform 1 0 122 0 1 9171
box -34 -63 34 63
use M2_M1431059130208_3v512x8m81  M2_M1431059130208_3v512x8m81_4
timestamp 1764525316
transform 1 0 281 0 1 11285
box -34 -63 34 63
use M2_M1431059130208_3v512x8m81  M2_M1431059130208_3v512x8m81_5
timestamp 1764525316
transform 1 0 276 0 1 8389
box -34 -63 34 63
use M2_M1431059130208_3v512x8m81  M2_M1431059130208_3v512x8m81_6
timestamp 1764525316
transform 1 0 430 0 1 9800
box -34 -63 34 63
use M2_M1431059130208_3v512x8m81  M2_M1431059130208_3v512x8m81_7
timestamp 1764525316
transform 1 0 281 0 1 10780
box -34 -63 34 63
use M2_M14310591302020_3v512x8m81  M2_M14310591302020_3v512x8m81_0
timestamp 1764525316
transform 1 0 285 0 1 4902
box -35 -56 35 55
use M2_M14310591302020_3v512x8m81  M2_M14310591302020_3v512x8m81_1
timestamp 1764525316
transform 1 0 280 0 1 5910
box -35 -56 35 55
use M2_M14310591302020_3v512x8m81  M2_M14310591302020_3v512x8m81_5
timestamp 1764525316
transform 0 -1 120 1 0 7459
box -35 -56 35 55
use M2_M14310591302020_3v512x8m81  M2_M14310591302020_3v512x8m81_6
timestamp 1764525316
transform 1 0 324 0 1 7183
box -35 -56 35 55
use M2_M14310591302020_3v512x8m81  M2_M14310591302020_3v512x8m81_9
timestamp 1764525316
transform 1 0 285 0 1 6993
box -35 -56 35 55
use M3_M2431059130201_3v512x8m81  M3_M2431059130201_3v512x8m81_1
timestamp 1764525316
transform 1 0 324 0 1 7190
box -35 -63 35 63
use nmos_1p2$$47119404_3v512x8m81  nmos_1p2$$47119404_3v512x8m81_1
timestamp 1764525316
transform 1 0 264 0 -1 6826
box -102 -44 130 679
use nmos_1p2$$47119404_3v512x8m81  nmos_1p2$$47119404_3v512x8m81_3
timestamp 1764525316
transform 1 0 264 0 -1 8190
box -102 -44 130 679
use nmos_5p0431059130202_3v512x8m81  nmos_5p0431059130202_3v512x8m81_0
timestamp 1764525316
transform 1 0 204 0 1 4329
box -124 -44 285 98
use pmos_1p2$$46889004_3v512x8m81  pmos_1p2$$46889004_3v512x8m81_1
timestamp 1764525316
transform 1 0 264 0 -1 5811
box -188 -86 216 721
use pmos_5p0431059130201_3v512x8m81  pmos_5p0431059130201_3v512x8m81_0
timestamp 1764525316
transform 1 0 248 0 -1 10077
box -174 -86 230 721
use pmos_5p0431059130201_3v512x8m81  pmos_5p0431059130201_3v512x8m81_1
timestamp 1764525316
transform 1 0 250 0 -1 9231
box -174 -86 230 721
use via1_2_3v512x8m81  via1_2_3v512x8m81_0
timestamp 1764525316
transform 1 0 174 0 1 4115
box 0 0 65 89
use via1_R90_3v512x8m81  via1_R90_3v512x8m81_0
timestamp 1764525316
transform -1 0 328 0 -1 6117
box 0 0 65 89
use via1_R90_3v512x8m81  via1_R90_3v512x8m81_2
timestamp 1764525316
transform 0 -1 343 1 0 11435
box 0 0 65 89
use via1_R90_3v512x8m81  via1_R90_3v512x8m81_3
timestamp 1764525316
transform 0 -1 343 1 0 11621
box 0 0 65 89
use via2_R90_3v512x8m81  via2_R90_3v512x8m81_0
timestamp 1764525316
transform 0 -1 333 1 0 11435
box 0 0 65 89
use via2_R90_3v512x8m81  via2_R90_3v512x8m81_1
timestamp 1764525316
transform 0 -1 333 1 0 11621
box 0 0 65 89
<< labels >>
rlabel metal1 s 229 10312 229 10312 4 pcb
port 8 nsew
rlabel metal3 s 318 11384 318 11384 4 vdd
port 2 nsew
rlabel metal2 s 125 11421 125 11421 4 bb
port 4 nsew
rlabel metal2 s 441 11421 441 11421 4 b
port 3 nsew
rlabel metal1 s 318 5007 318 5007 4 vdd
port 2 nsew
rlabel metal2 s 261 4923 261 4923 4 ypass
port 6 nsew
rlabel metal2 s 54 4251 54 4251 4 db
port 5 nsew
rlabel metal2 s 44 4251 44 4251 6 db
port 5 nsew
rlabel metal3 s 352 7303 352 7303 4 vss
port 1 nsew
rlabel metal3 -6 4244 -6 4245 0 vss
port 1 nsew
<< properties >>
string path 0.000 27.385 0.000 -0.005 
<< end >>
