magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal1 >>
rect -44 1321 45 1341
rect -44 -1321 -26 1321
rect 26 -1321 45 1321
rect -44 -1341 45 -1321
<< via1 >>
rect -26 -1321 26 1321
<< metal2 >>
rect -44 1321 45 1341
rect -44 -1321 -26 1321
rect 26 -1321 45 1321
rect -44 -1341 45 -1321
<< end >>
