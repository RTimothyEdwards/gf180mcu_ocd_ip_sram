magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal1 >>
rect -113 408 113 417
rect -113 -408 -105 408
rect 105 -408 113 408
rect -113 -417 113 -408
<< via1 >>
rect -105 -408 105 408
<< metal2 >>
rect -113 408 113 417
rect -113 -408 -105 408
rect 105 -408 113 408
rect -113 -417 113 -408
<< end >>
