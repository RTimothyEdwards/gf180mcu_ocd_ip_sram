magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< polysilicon >>
rect -240 23 240 46
rect -240 -23 -194 23
rect 194 -23 240 23
rect -240 -46 240 -23
<< polycontact >>
rect -194 -23 194 23
<< metal1 >>
rect -213 23 213 40
rect -213 -23 -194 23
rect 194 -23 213 23
rect -213 -39 213 -23
<< end >>
