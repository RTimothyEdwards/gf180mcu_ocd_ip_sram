magic
tech gf180mcuD
magscale 1 10
timestamp 1763477050
<< metal2 >>
rect -5 1821 151 4266
rect 346 2590 503 5538
rect 707 1821 864 4263
use M2_M14310591302097_512x8m81  M2_M14310591302097_512x8m81_0
timestamp 1763476864
transform 1 0 784 0 1 2162
box -70 -330 70 330
use M2_M14310591302097_512x8m81  M2_M14310591302097_512x8m81_1
timestamp 1763476864
transform 1 0 72 0 1 2162
box -70 -330 70 330
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_0
timestamp 1763476864
transform 1 0 424 0 1 4630
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_1
timestamp 1763476864
transform 1 0 786 0 1 3500
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_2
timestamp 1763476864
transform 1 0 74 0 1 3500
box -70 -113 70 113
use M3_M24310591302096_512x8m81  M3_M24310591302096_512x8m81_0
timestamp 1763476864
transform 1 0 424 0 1 2886
box -70 -287 70 287
<< properties >>
string path 5.615 28.025 5.615 10.575 
<< end >>
