magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< metal1 >>
rect -1815 247 1815 275
rect -1815 -247 -1789 247
rect 1789 -247 1815 247
rect -1815 -275 1815 -247
<< via1 >>
rect -1789 -247 1789 247
<< metal2 >>
rect -1815 247 1815 275
rect -1815 -247 -1789 247
rect 1789 -247 1815 247
rect -1815 -275 1815 -247
<< end >>
