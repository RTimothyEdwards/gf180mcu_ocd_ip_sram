magic
tech gf180mcuD
magscale 1 10
timestamp 1766784746
<< nwell >>
rect -161 5039 54 8484
rect -121 2318 3694 2520
rect -121 1751 3715 2318
rect -121 1473 739 1751
rect 902 1503 3715 1751
rect 902 1473 3694 1503
rect -121 1104 3694 1473
<< metal1 >>
rect -16 6908 3476 6960
<< metal2 >>
rect 7 8278 63 8338
rect 340 8278 396 8338
rect 464 8278 520 8338
rect 797 8278 853 8338
rect 909 8278 965 8338
rect 1242 8278 1298 8338
rect 1366 8278 1422 8338
rect 1699 8278 1755 8338
rect 1811 8278 1867 8338
rect 2144 8278 2200 8338
rect 2268 8278 2324 8338
rect 2601 8278 2657 8338
rect 2713 8278 2769 8338
rect 3046 8278 3102 8338
rect 3158 8278 3214 8338
rect 3528 8278 3584 8338
rect 40 3516 103 3576
rect 757 3516 820 3576
rect 942 3516 1005 3576
rect 1659 3516 1722 3576
rect 1844 3516 1907 3576
rect 2561 3516 2624 3576
rect 2746 3516 2809 3576
rect 3501 3519 3564 3579
rect 774 1499 845 1710
rect 1689 1495 1750 1707
rect 2591 1495 2652 1699
<< metal3 >>
rect -575 5420 4956 5618
use M1_NACTIVE4310591302028_3v256x8m81  M1_NACTIVE4310591302028_3v256x8m81_0
timestamp 1765833244
transform 1 0 426 0 1 5519
box -122 -181 122 181
use M1_NACTIVE4310591302028_3v256x8m81  M1_NACTIVE4310591302028_3v256x8m81_1
timestamp 1765833244
transform 1 0 1332 0 1 5519
box -122 -181 122 181
use M1_NACTIVE4310591302028_3v256x8m81  M1_NACTIVE4310591302028_3v256x8m81_2
timestamp 1765833244
transform 1 0 2236 0 1 5519
box -122 -181 122 181
use M1_NACTIVE4310591302028_3v256x8m81  M1_NACTIVE4310591302028_3v256x8m81_3
timestamp 1765833244
transform 1 0 3140 0 1 5519
box -122 -181 122 181
use M2_M14310591302018_3v256x8m81  M2_M14310591302018_3v256x8m81_0
timestamp 1765833244
transform 1 0 426 0 1 5519
box -34 -99 34 99
use M2_M14310591302018_3v256x8m81  M2_M14310591302018_3v256x8m81_1
timestamp 1765833244
transform 1 0 1332 0 1 5519
box -34 -99 34 99
use M2_M14310591302018_3v256x8m81  M2_M14310591302018_3v256x8m81_2
timestamp 1765833244
transform 1 0 2236 0 1 5519
box -34 -99 34 99
use M2_M14310591302018_3v256x8m81  M2_M14310591302018_3v256x8m81_3
timestamp 1765833244
transform 1 0 3140 0 1 5519
box -34 -99 34 99
use M2_M14310591302020_3v256x8m81  M2_M14310591302020_3v256x8m81_0
timestamp 1765833244
transform 1 0 809 0 1 1648
box -35 -56 35 55
use M2_M14310591302020_3v256x8m81  M2_M14310591302020_3v256x8m81_2
timestamp 1765833244
transform 1 0 1719 0 1 1648
box -35 -56 35 55
use M2_M14310591302020_3v256x8m81  M2_M14310591302020_3v256x8m81_4
timestamp 1765833244
transform 1 0 2621 0 1 1648
box -35 -56 35 55
use M3_M2431059130201_3v256x8m81  M3_M2431059130201_3v256x8m81_0
timestamp 1765833244
transform 1 0 809 0 1 1581
box -35 -63 35 63
use M3_M2431059130201_3v256x8m81  M3_M2431059130201_3v256x8m81_1
timestamp 1765833244
transform 1 0 1719 0 1 1581
box -35 -63 35 63
use M3_M2431059130201_3v256x8m81  M3_M2431059130201_3v256x8m81_3
timestamp 1765833244
transform 1 0 2621 0 1 1581
box -35 -63 35 63
use M3_M24310591302029_3v256x8m81  M3_M24310591302029_3v256x8m81_0
timestamp 1765833244
transform 1 0 426 0 1 5519
box -35 -99 35 99
use M3_M24310591302029_3v256x8m81  M3_M24310591302029_3v256x8m81_1
timestamp 1765833244
transform 1 0 1332 0 1 5519
box -35 -99 35 99
use M3_M24310591302029_3v256x8m81  M3_M24310591302029_3v256x8m81_2
timestamp 1765833244
transform 1 0 2236 0 1 5519
box -35 -99 35 99
use M3_M24310591302029_3v256x8m81  M3_M24310591302029_3v256x8m81_3
timestamp 1765833244
transform 1 0 3140 0 1 5519
box -35 -99 35 99
use ypass_gate_3v256x8m81  ypass_gate_3v256x8m81_1
timestamp 1766784746
transform -1 0 3190 0 1 -3377
box -130 4011 633 11861
use ypass_gate_3v256x8m81  ypass_gate_3v256x8m81_2
timestamp 1766784746
transform -1 0 2288 0 1 -3377
box -130 4011 633 11861
use ypass_gate_3v256x8m81  ypass_gate_3v256x8m81_3
timestamp 1766784746
transform -1 0 1386 0 1 -3377
box -130 4011 633 11861
use ypass_gate_3v256x8m81  ypass_gate_3v256x8m81_4
timestamp 1766784746
transform 1 0 2180 0 1 -3377
box -130 4011 633 11861
use ypass_gate_3v256x8m81  ypass_gate_3v256x8m81_5
timestamp 1766784746
transform 1 0 1278 0 1 -3377
box -130 4011 633 11861
use ypass_gate_3v256x8m81  ypass_gate_3v256x8m81_6
timestamp 1766784746
transform 1 0 376 0 1 -3377
box -130 4011 633 11861
use ypass_gate_3v256x8m81  ypass_gate_3v256x8m81_7
timestamp 1766784746
transform -1 0 484 0 1 -3377
box -130 4011 633 11861
use ypass_gate_a_3v256x8m81  ypass_gate_a_3v256x8m81_0
timestamp 1765900146
transform 1 0 3090 0 1 -3377
box -130 4017 627 11860
<< labels >>
rlabel metal2 70 3546 70 3546 0 ypass[0]
rlabel metal2 788 3543 788 3543 0 ypass[1]
rlabel metal2 973 3543 973 3543 0 ypass[2]
rlabel metal2 1689 3544 1689 3544 0 ypass[3]
rlabel metal2 1874 3544 1874 3544 0 ypass[4]
rlabel metal2 2591 3543 2591 3543 0 ypass[5]
rlabel metal2 2776 3543 2776 3543 0 ypass[6]
rlabel metal2 3533 3546 3533 3546 0 ypass[7]
rlabel metal2 33 8307 33 8307 0 b[0]
rlabel metal2 366 8306 366 8306 0 bb[0]
rlabel metal2 490 8307 490 8307 0 bb[1]
rlabel metal2 824 8306 824 8306 0 b[1]
rlabel metal2 935 8307 935 8307 0 b[2]
rlabel metal2 1271 8306 1271 8306 0 bb[2]
rlabel metal2 1393 8306 1393 8306 0 bb[3]
rlabel metal2 1728 8305 1728 8305 0 b[3]
rlabel metal2 1838 8306 1838 8306 0 b[4]
rlabel metal2 2171 8306 2171 8306 0 bb[4]
rlabel metal2 2294 8306 2294 8306 0 bb[5]
rlabel metal2 2629 8305 2629 8305 0 b[5]
rlabel metal2 2740 8305 2740 8305 0 b[6]
rlabel metal2 3073 8306 3073 8306 0 bb[6]
rlabel metal2 3186 8306 3186 8306 0 bb[7]
rlabel metal2 3554 8307 3554 8307 0 b[7]
<< end >>
