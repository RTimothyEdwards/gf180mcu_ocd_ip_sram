magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< error_s >>
rect -89 0 -43 89
rect 71 0 117 89
<< polysilicon >>
rect -14 89 41 123
rect -14 -34 41 0
use nmos_5p0431059130208_3v512x8m81  nmos_5p0431059130208_3v512x8m81_0
timestamp 1764525316
transform 1 0 -14 0 1 0
box -88 -44 144 133
<< end >>
