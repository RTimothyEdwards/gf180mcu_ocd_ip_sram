magic
tech gf180mcuD
magscale 1 10
timestamp 1763588843
<< error_s >>
rect 16287 15009 16298 15012
rect 16343 14647 16354 15009
rect 1572 14114 1611 14115
rect 1645 14114 1684 14115
rect 1770 14114 1809 14115
rect 1843 14114 1882 14115
rect 1968 14114 2007 14115
rect 2041 14114 2080 14115
rect 2852 14114 2891 14115
rect 2925 14114 2964 14115
rect 3050 14114 3089 14115
rect 3123 14114 3162 14115
rect 3248 14114 3287 14115
rect 3321 14114 3360 14115
rect 6737 14114 6776 14115
rect 6810 14114 6849 14115
rect 6935 14114 6974 14115
rect 7008 14114 7047 14115
rect 7133 14114 7172 14115
rect 7206 14114 7245 14115
rect 8017 14114 8056 14115
rect 8090 14114 8129 14115
rect 8215 14114 8254 14115
rect 8288 14114 8327 14115
rect 8413 14114 8452 14115
rect 8486 14114 8525 14115
<< nwell >>
rect 17442 19330 18301 19778
rect 17262 8699 17293 8720
rect 18106 8699 18193 8720
rect 18983 8699 19055 8720
rect 14494 7349 15036 7710
rect 16382 7653 19055 8699
rect 14517 6396 14632 6429
rect 17262 5806 17293 7653
rect 18106 5377 18193 7653
rect 18983 5471 19055 7653
rect 5846 2204 6015 2612
<< metal1 >>
rect 282 2508 375 20398
rect 1143 20257 1270 20304
rect 4808 14067 4899 14208
rect 535 13973 4899 14067
rect 535 9206 625 13973
rect 6001 13908 6092 14199
rect 704 13814 6092 13908
rect 704 9470 795 13814
rect 9952 13749 10042 14187
rect 873 13656 10042 13749
rect 11136 13793 11226 14241
rect 17292 13952 17383 14450
rect 18476 14111 18566 14439
rect 19660 14269 19753 14472
rect 19660 14176 20202 14269
rect 18476 14017 20033 14111
rect 17292 13859 19864 13952
rect 11136 13700 19695 13793
rect 873 9675 963 13656
rect 873 9586 1290 9675
rect 704 9361 1121 9470
rect 535 9099 952 9206
rect 861 2264 952 9099
rect 1031 2264 1121 9361
rect 1199 2264 1290 9586
rect 14693 8441 14743 8570
rect 15017 8441 15068 8575
rect 15336 8441 15386 8561
rect 14693 8391 15386 8441
rect 14710 8390 15369 8391
rect 15701 2862 15748 2864
rect 14532 2813 15748 2862
rect 9200 1985 10308 2033
rect 15701 2007 15748 2813
rect 19604 2121 19695 13700
rect 19773 2121 19864 13859
rect 19943 2121 20033 14017
rect 20111 2121 20202 14176
rect 20664 2508 20757 20366
rect 282 1612 6454 1931
rect 9200 648 9248 1985
rect 19488 1612 20590 1931
<< metal2 >>
rect 451 2667 1043 21087
rect 12009 20205 12100 20298
rect 12255 20205 12345 20298
rect 13153 20205 13244 20298
rect 13402 20205 13492 20298
rect 14298 20205 14389 20298
rect 14538 20205 14628 20298
rect 15439 20205 15529 20298
rect 15691 20205 15781 20298
rect 1635 20046 1725 20140
rect 1883 20046 1974 20140
rect 2887 20046 2978 20140
rect 3141 20046 3231 20140
rect 6799 20046 6890 20140
rect 7049 20046 7139 20140
rect 8052 20046 8143 20140
rect 8306 20046 8397 20140
rect 282 702 375 2509
rect 451 1612 760 2667
rect 861 702 952 2509
rect 1031 702 1121 2509
rect 1199 702 1290 2509
rect 2359 702 2452 3052
rect 3542 702 3636 3068
rect 4727 702 4821 3059
rect 6274 2924 6364 3076
rect 5693 2830 6364 2924
rect 11423 2855 11480 2857
rect 5693 1008 5783 2830
rect 11353 2816 11480 2855
rect 6216 1816 6454 2724
rect 11423 744 11480 2816
rect 15128 1600 15375 4119
rect 19972 2667 20588 21087
rect 15998 702 16092 2132
rect 19604 702 19695 2519
rect 19773 702 19864 2519
rect 19943 702 20033 2519
rect 20111 702 20202 2519
rect 20279 1612 20588 2667
rect 20664 820 20757 2509
<< metal3 >>
rect 451 20451 20588 21087
rect 282 20324 20757 20366
rect 282 20150 20667 20324
rect 20753 20150 20757 20324
rect 19677 12097 19767 12190
rect 19677 11859 19767 11952
rect 19677 11621 19767 11714
rect 19677 11383 19767 11476
rect 19677 11145 19767 11238
rect 19677 10907 19767 11000
rect 19677 10668 19767 10762
rect 19677 10430 19767 10524
use gen_256x8_256x8m81  gen_256x8_256x8m81_0
timestamp 1763588843
transform 1 0 9916 0 1 2199
box -12453 -1374 12336 11499
use M1_NACTIVE4310591302047_256x8m81  M1_NACTIVE4310591302047_256x8m81_0
timestamp 1763564386
transform 0 -1 18221 1 0 19550
box -62 -36 62 36
use M1_NACTIVE4310591302047_256x8m81  M1_NACTIVE4310591302047_256x8m81_1
timestamp 1763564386
transform 0 -1 17500 1 0 19559
box -62 -36 62 36
use M1_PACTIVE4310591302048_256x8m81  M1_PACTIVE4310591302048_256x8m81_0
timestamp 1763565688
transform 1 0 2440 0 1 20281
box -1152 -36 1153 36
use M1_PACTIVE4310591302048_256x8m81  M1_PACTIVE4310591302048_256x8m81_1
timestamp 1763565688
transform 1 0 7592 0 1 20281
box -1152 -36 1153 36
use M1_PACTIVE4310591302049_256x8m81  M1_PACTIVE4310591302049_256x8m81_0
timestamp 1763564386
transform 1 0 16713 0 1 20268
box -457 -36 457 36
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_0
timestamp 1763564386
transform -1 0 20710 0 1 20272
box -43 -122 43 122
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_1
timestamp 1763564386
transform -1 0 20710 0 1 2387
box -43 -122 43 122
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_2
timestamp 1763564386
transform 1 0 329 0 1 20262
box -43 -122 43 122
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_3
timestamp 1763564386
transform 1 0 329 0 1 2387
box -43 -122 43 122
use M2_M1$$199746604_256x8m81  M2_M1$$199746604_256x8m81_0
timestamp 1763564386
transform 1 0 605 0 1 1771
box -119 -123 119 123
use M2_M1$$199746604_256x8m81  M2_M1$$199746604_256x8m81_1
timestamp 1763564386
transform 1 0 20433 0 1 1771
box -119 -123 119 123
use M2_M1$$199746604_256x8m81  M2_M1$$199746604_256x8m81_2
timestamp 1763564386
transform 1 0 6335 0 1 1697
box -119 -123 119 123
use M2_M1$$201262124_256x8m81  M2_M1$$201262124_256x8m81_0
timestamp 1763564386
transform 1 0 6335 0 1 1884
box -119 -46 119 46
use M2_M1$$202405932_256x8m81  M2_M1$$202405932_256x8m81_0
timestamp 1763564386
transform 1 0 20157 0 1 2320
box -44 -198 44 198
use M2_M1$$202405932_256x8m81  M2_M1$$202405932_256x8m81_1
timestamp 1763564386
transform 1 0 19988 0 1 2320
box -44 -198 44 198
use M2_M1$$202405932_256x8m81  M2_M1$$202405932_256x8m81_2
timestamp 1763564386
transform 1 0 19819 0 1 2320
box -44 -198 44 198
use M2_M1$$202405932_256x8m81  M2_M1$$202405932_256x8m81_3
timestamp 1763564386
transform 1 0 19649 0 1 2320
box -44 -198 44 198
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_0
timestamp 1763564386
transform 1 0 1245 0 1 2387
box -45 -122 45 123
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_1
timestamp 1763564386
transform 1 0 1075 0 1 2387
box -45 -122 45 123
use M2_M1$$202406956_256x8m81  M2_M1$$202406956_256x8m81_2
timestamp 1763564386
transform 1 0 907 0 1 2387
box -45 -122 45 123
use M3_M2$$43368492_256x8m81  M3_M2$$43368492_256x8m81_0
timestamp 1763564386
transform -1 0 20710 0 1 20272
box -44 -123 44 123
use M3_M2$$43368492_256x8m81  M3_M2$$43368492_256x8m81_1
timestamp 1763564386
transform 1 0 329 0 1 20272
box -44 -123 44 123
use M3_M2$$201255980_256x8m81  M3_M2$$201255980_256x8m81_0
timestamp 1763564386
transform -1 0 20640 0 1 1028
box -119 -46 119 46
use M3_M2$$201255980_256x8m81  M3_M2$$201255980_256x8m81_1
timestamp 1763564386
transform 1 0 399 0 1 1028
box -119 -46 119 46
use M3_M2$$201255980_256x8m81  M3_M2$$201255980_256x8m81_2
timestamp 1763564386
transform 1 0 5738 0 1 1028
box -119 -46 119 46
use M3_M2$$201401388_256x8m81  M3_M2$$201401388_256x8m81_0
timestamp 1763564386
transform 1 0 20280 0 1 20769
box -266 -275 266 275
use M3_M2$$201401388_256x8m81  M3_M2$$201401388_256x8m81_1
timestamp 1763564386
transform 1 0 759 0 1 20769
box -266 -275 266 275
use M3_M2$$201401388_256x8m81  M3_M2$$201401388_256x8m81_2
timestamp 1763564386
transform 1 0 20280 0 1 8482
box -266 -275 266 275
use M3_M24310591302050_256x8m81  M3_M24310591302050_256x8m81_0
timestamp 1763564386
transform 1 0 15254 0 1 1756
box -99 -99 99 99
use M3_M24310591302050_256x8m81  M3_M24310591302050_256x8m81_1
timestamp 1763564386
transform 1 0 15254 0 1 2372
box -99 -99 99 99
use prexdec_top_256x8m81  prexdec_top_256x8m81_0
timestamp 1763587904
transform 1 0 949 0 1 12306
box 21 1806 19120 8780
use ypredec1_256x8m81  ypredec1_256x8m81_0
timestamp 1763578215
transform 1 0 1092 0 1 2092
box 125 53 18674 11572
<< labels >>
rlabel metal3 s 1263 8767 1263 8767 4 LYS[0]
port 11 nsew
rlabel metal3 s 1263 9005 1263 9005 4 LYS[1]
port 12 nsew
rlabel metal3 s 1263 9243 1263 9243 4 LYS[2]
port 13 nsew
rlabel metal3 s 1263 9481 1263 9481 4 LYS[3]
port 14 nsew
rlabel metal3 s 1263 10195 1263 10195 4 LYS[6]
port 15 nsew
rlabel metal3 s 1263 9957 1263 9957 4 LYS[5]
port 16 nsew
rlabel metal3 s 1263 9719 1263 9719 4 LYS[4]
port 17 nsew
rlabel metal3 s 18802 20769 18802 20769 4 men
port 18 nsew
rlabel metal3 s 1263 10434 1263 10434 4 LYS[7]
port 19 nsew
flabel metal3 s 4365 13286 4365 13286 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 4365 16804 4365 16804 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 4365 19672 4365 19672 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 4365 18246 4365 18246 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 4365 11179 4365 11179 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 4365 18978 4365 18978 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 4365 14201 4365 14201 0 FreeSans 313 0 0 0 VSS
port 1 nsew
rlabel metal2 s 6808 20123 6808 20123 4 xb[3]
port 22 nsew
rlabel metal2 s 7114 20128 7114 20128 4 xb[2]
port 23 nsew
rlabel metal2 s 8376 20111 8376 20111 4 xb[0]
port 24 nsew
rlabel metal2 s 12054 20251 12054 20251 4 xa[7]
port 25 nsew
rlabel metal2 s 12300 20251 12300 20251 4 xa[6]
port 26 nsew
rlabel metal2 s 13198 20251 13198 20251 4 xa[5]
port 27 nsew
rlabel metal2 s 13447 20251 13447 20251 4 xa[4]
port 28 nsew
rlabel metal2 s 14343 20251 14343 20251 4 xa[3]
port 29 nsew
rlabel metal2 s 14583 20251 14583 20251 4 xa[2]
port 30 nsew
rlabel metal2 s 8068 20098 8068 20098 4 xb[1]
port 33 nsew
rlabel metal2 s 7094 20093 7094 20093 4 xb[2]
port 23 nsew
rlabel metal2 s 8351 20090 8351 20090 4 xb[0]
port 24 nsew
rlabel metal2 s 1680 20093 1680 20093 4 xc[3]
port 34 nsew
rlabel metal2 s 2933 20090 2933 20090 4 xc[1]
port 35 nsew
rlabel metal2 s 1929 20093 1929 20093 4 xc[2]
port 36 nsew
rlabel metal2 s 3186 20090 3186 20090 4 xc[0]
port 37 nsew
rlabel metal2 s 15736 20251 15736 20251 4 xa[0]
port 38 nsew
rlabel metal2 s 15484 20251 15484 20251 4 xa[1]
port 39 nsew
rlabel metal2 s 8098 20090 8098 20090 4 xb[1]
port 33 nsew
rlabel metal2 s 6845 20093 6845 20093 4 xb[3]
port 22 nsew
flabel metal3 s 4365 14442 4365 14442 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal1 s 9219 762 9219 762 0 FreeSans 700 0 0 0 GWEN
port 51 nsew
flabel metal1 s 15717 2437 15717 2437 0 FreeSans 700 0 0 0 GWE
port 50 nsew
rlabel metal2 s 1075 748 1075 748 4 A[8]
port 49 nsew
rlabel metal2 s 19819 748 19819 748 4 A[5]
port 48 nsew
rlabel metal2 s 19988 748 19988 748 4 A[4]
port 47 nsew
rlabel metal2 s 20157 748 20157 748 4 A[3]
port 46 nsew
rlabel metal2 s 19649 748 19649 748 4 A[6]
port 45 nsew
rlabel metal2 s 3589 748 3589 748 4 A[1]
port 44 nsew
rlabel metal2 s 2405 748 2405 748 4 A[2]
port 43 nsew
rlabel metal2 s 329 748 329 748 4 CLK
port 42 nsew
rlabel metal2 s 1245 748 1245 748 4 A[7]
port 41 nsew
rlabel metal2 s 907 748 907 748 4 A[9]
port 40 nsew
rlabel metal2 s 16046 748 16046 748 4 CEN
port 32 nsew
rlabel metal2 s 4774 748 4774 748 4 A[0]
port 31 nsew
flabel metal2 s 11449 762 11449 762 0 FreeSans 700 0 0 0 IGWEN
port 21 nsew
flabel metal3 s 4365 6277 4365 6277 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 4365 3413 4365 3413 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 5796 2441 5796 2441 0 FreeSans 313 0 0 0 VDD
port 2 nsew
flabel metal3 s 4365 2676 4365 2676 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 4365 4149 4365 4149 0 FreeSans 313 0 0 0 VSS
port 1 nsew
flabel metal3 s 4365 8014 4365 8014 0 FreeSans 313 0 0 0 VSS
port 1 nsew
rlabel metal3 s 19569 5213 19569 5213 4 tblhl
port 20 nsew
flabel metal3 s 5796 1454 5796 1454 0 FreeSans 313 0 0 0 VDD
port 2 nsew
rlabel metal3 s 19722 12144 19722 12144 4 RYS[7]
port 3 nsew
rlabel metal3 s 19722 11905 19722 11905 4 RYS[6]
port 4 nsew
rlabel metal3 s 19722 11667 19722 11667 4 RYS[5]
port 5 nsew
rlabel metal3 s 19722 11429 19722 11429 4 RYS[4]
port 6 nsew
rlabel metal3 s 19722 11191 19722 11191 4 RYS[3]
port 7 nsew
rlabel metal3 s 19722 10953 19722 10953 4 RYS[2]
port 8 nsew
rlabel metal3 s 19722 10715 19722 10715 4 RYS[1]
port 9 nsew
rlabel metal3 s 19722 10477 19722 10477 4 RYS[0]
port 10 nsew
flabel metal3 s 5488 1266 5488 1266 0 FreeSans 313 0 0 0 VSS
port 1 nsew
<< properties >>
string path 81.095 8.115 81.735 8.115 81.735 -9.165 
<< end >>
