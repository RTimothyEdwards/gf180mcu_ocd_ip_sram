magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nwell >>
rect -426 338 1350 339
rect -426 337 1374 338
rect -426 335 1398 337
rect -426 -86 1422 335
<< pmos >>
rect -252 0 -196 253
rect -92 0 -36 253
rect 69 0 125 253
rect 229 0 285 253
rect 390 0 446 253
rect 550 0 606 253
rect 711 0 767 253
rect 871 0 927 253
rect 1032 0 1088 253
rect 1192 0 1248 253
<< pdiff >>
rect -340 240 -252 253
rect -340 13 -327 240
rect -281 13 -252 240
rect -340 0 -252 13
rect -196 240 -92 253
rect -196 13 -167 240
rect -121 13 -92 240
rect -196 0 -92 13
rect -36 240 69 253
rect -36 13 -7 240
rect 39 13 69 240
rect -36 0 69 13
rect 125 240 229 253
rect 125 13 154 240
rect 200 13 229 240
rect 125 0 229 13
rect 285 240 390 253
rect 285 13 314 240
rect 360 13 390 240
rect 285 0 390 13
rect 446 240 550 253
rect 446 13 475 240
rect 521 13 550 240
rect 446 0 550 13
rect 606 240 711 253
rect 606 13 635 240
rect 681 13 711 240
rect 606 0 711 13
rect 767 240 871 253
rect 767 13 796 240
rect 842 13 871 240
rect 767 0 871 13
rect 927 240 1032 253
rect 927 13 956 240
rect 1002 13 1032 240
rect 927 0 1032 13
rect 1088 240 1192 253
rect 1088 13 1117 240
rect 1163 13 1192 240
rect 1088 0 1192 13
rect 1248 240 1336 253
rect 1248 13 1277 240
rect 1323 13 1336 240
rect 1248 0 1336 13
<< pdiffc >>
rect -327 13 -281 240
rect -167 13 -121 240
rect -7 13 39 240
rect 154 13 200 240
rect 314 13 360 240
rect 475 13 521 240
rect 635 13 681 240
rect 796 13 842 240
rect 956 13 1002 240
rect 1117 13 1163 240
rect 1277 13 1323 240
<< polysilicon >>
rect -252 253 -196 297
rect -92 253 -36 297
rect 69 253 125 297
rect 229 253 285 297
rect 390 253 446 297
rect 550 253 606 297
rect 711 253 767 297
rect 871 253 927 297
rect 1032 253 1088 297
rect 1192 253 1248 297
rect -252 -45 -196 0
rect -92 -45 -36 0
rect 69 -45 125 0
rect 229 -45 285 0
rect 390 -45 446 0
rect 550 -45 606 0
rect 711 -45 767 0
rect 871 -45 927 0
rect 1032 -45 1088 0
rect 1192 -45 1248 0
<< metal1 >>
rect -327 240 -281 253
rect -327 0 -281 13
rect -167 240 -121 253
rect -167 0 -121 13
rect -7 240 39 253
rect -7 0 39 13
rect 154 240 200 253
rect 154 0 200 13
rect 314 240 360 253
rect 314 0 360 13
rect 475 240 521 253
rect 475 0 521 13
rect 635 240 681 253
rect 635 0 681 13
rect 796 240 842 253
rect 796 0 842 13
rect 956 240 1002 253
rect 956 0 1002 13
rect 1117 240 1163 253
rect 1117 0 1163 13
rect 1277 240 1323 253
rect 1277 0 1323 13
<< labels >>
flabel pdiffc 498 126 498 126 0 FreeSans 186 0 0 0 D
flabel pdiffc 349 126 349 126 0 FreeSans 186 0 0 0 S
flabel pdiffc 189 126 189 126 0 FreeSans 186 0 0 0 D
flabel pdiffc 28 126 28 126 0 FreeSans 186 0 0 0 S
flabel pdiffc -132 126 -132 126 0 FreeSans 186 0 0 0 D
flabel pdiffc -292 126 -292 126 0 FreeSans 186 0 0 0 S
flabel pdiffc 807 126 807 126 0 FreeSans 186 0 0 0 D
flabel pdiffc 1128 126 1128 126 0 FreeSans 186 0 0 0 D
flabel pdiffc 1289 126 1289 126 0 FreeSans 186 0 0 0 S
flabel pdiffc 645 126 645 126 0 FreeSans 186 0 0 0 S
flabel pdiffc 967 126 967 126 0 FreeSans 186 0 0 0 S
<< end >>
