magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< nwell >>
rect -137 -63 165 678
<< polysilicon >>
rect -14 615 41 648
rect -14 -33 41 0
use pmos_5p043105913020101_256x8m81  pmos_5p043105913020101_256x8m81_0
timestamp 1763564386
transform 1 0 -14 0 1 0
box -174 -86 230 701
<< end >>
