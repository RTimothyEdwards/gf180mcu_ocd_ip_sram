magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal1 >>
rect -123 40 122 45
rect -123 26 123 40
rect -123 -26 -102 26
rect 102 -26 123 26
rect -123 -40 123 -26
rect -123 -45 122 -40
<< via1 >>
rect -102 -26 102 26
<< metal2 >>
rect -123 26 122 45
rect -123 -26 -102 26
rect 102 -26 122 26
rect -123 -45 122 -26
<< end >>
