magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< error_s >>
rect 390 948 420 1068
rect 389 724 420 948
rect 389 115 420 129
<< polysilicon >>
rect 533 4126 589 5015
rect 893 4126 949 5015
<< metal1 >>
rect 227 5055 529 5964
rect 605 4993 686 5098
rect 605 4909 901 4993
rect 245 2573 529 4846
rect 605 3969 686 4909
rect 965 3998 1045 5098
rect -74 2436 1276 2501
rect -74 2295 1276 2360
rect -74 2154 1276 2219
rect -74 2013 1276 2078
rect -74 1871 1276 1936
rect -74 1730 1276 1795
<< metal2 >>
rect 294 5302 529 5853
rect 294 951 385 4998
rect 800 989 890 2657
rect 1143 1130 1233 2839
rect 800 896 1233 989
<< metal3 >>
rect 0 5263 1276 5898
rect 0 3120 1184 5026
rect 4 2821 1233 2914
rect 9 2564 1270 2657
rect 800 2563 890 2564
use alatch_512x8m81  alatch_512x8m81_0
timestamp 1763476864
transform 1 0 49 0 1 -442
box -63 0 1196 2077
use M1_NWELL10_512x8m81  M1_NWELL10_512x8m81_0
timestamp 1763476864
transform 1 0 233 0 1 3599
box -154 -1130 154 1130
use M1_POLY2$$46559276_512x8m81  M1_POLY2$$46559276_512x8m81_0
timestamp 1763476864
transform 1 0 805 0 1 4951
box -123 -48 123 48
use M1_POLY2$$46559276_512x8m81  M1_POLY2$$46559276_512x8m81_1
timestamp 1763476864
transform 1 0 448 0 1 4951
box -123 -48 123 48
use M1_PSUB$$47335468_512x8m81  M1_PSUB$$47335468_512x8m81_0
timestamp 1763476864
transform 1 0 276 0 1 5537
box -55 -400 56 400
use M2_M1$$34864172_512x8m81  M2_M1$$34864172_512x8m81_0
timestamp 1763476864
transform 1 0 413 0 1 4951
box -119 -46 119 46
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1763476864
transform 1 0 339 0 1 1042
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_1
timestamp 1763476864
transform 1 0 645 0 1 2696
box -43 -122 43 122
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_2
timestamp 1763476864
transform 1 0 1005 0 1 2696
box -43 -122 43 122
use M2_M1$$43377708_512x8m81  M2_M1$$43377708_512x8m81_0
timestamp 1763476864
transform 1 0 853 0 1 4349
box -44 -427 44 427
use M2_M1$$43377708_512x8m81  M2_M1$$43377708_512x8m81_1
timestamp 1763476864
transform 1 0 493 0 1 4349
box -44 -427 44 427
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_0
timestamp 1763476864
transform 1 0 339 0 1 5578
box -44 -275 44 275
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_1
timestamp 1763476864
transform 1 0 484 0 1 5578
box -44 -275 44 275
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_2
timestamp 1763476864
transform 1 0 848 0 1 5578
box -44 -275 44 275
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_0
timestamp 1763476864
transform 1 0 1188 0 1 2867
box -44 -123 44 123
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_1
timestamp 1763476864
transform 1 0 845 0 1 2534
box -44 -123 44 123
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_0
timestamp 1763476864
transform 1 0 339 0 1 5578
box -45 -275 45 275
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_1
timestamp 1763476864
transform 1 0 484 0 1 5578
box -45 -275 45 275
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_2
timestamp 1763476864
transform 1 0 848 0 1 5578
box -45 -275 45 275
use M3_M2$$47334444_512x8m81  M3_M2$$47334444_512x8m81_0
timestamp 1763476864
transform 1 0 853 0 1 4349
box -45 -427 45 427
use M3_M2$$47334444_512x8m81  M3_M2$$47334444_512x8m81_1
timestamp 1763476864
transform 1 0 493 0 1 4349
box -45 -427 45 427
use nmos_1p2$$47336492_512x8m81  nmos_1p2$$47336492_512x8m81_0
timestamp 1763476864
transform 1 0 907 0 1 5049
box -102 -44 130 658
use nmos_1p2$$47336492_512x8m81  nmos_1p2$$47336492_512x8m81_1
timestamp 1763476864
transform 1 0 547 0 1 5049
box -102 -44 130 658
use pmos_1p2$$47337516_512x8m81  pmos_1p2$$47337516_512x8m81_0
timestamp 1763476864
transform 1 0 907 0 1 2567
box -188 -86 216 1610
use pmos_1p2$$47337516_512x8m81  pmos_1p2$$47337516_512x8m81_1
timestamp 1763476864
transform 1 0 547 0 1 2567
box -188 -86 216 1610
<< end >>
