magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< nwell >>
rect -314 -86 892 297
<< pmos >>
rect -140 0 -84 211
rect 20 0 76 211
rect 181 0 237 211
rect 341 0 397 211
rect 502 0 558 211
rect 662 0 718 211
<< pdiff >>
rect -228 198 -140 211
rect -228 14 -215 198
rect -169 14 -140 198
rect -228 0 -140 14
rect -84 198 20 211
rect -84 14 -55 198
rect -9 14 20 198
rect -84 0 20 14
rect 76 198 181 211
rect 76 14 105 198
rect 151 14 181 198
rect 76 0 181 14
rect 237 198 341 211
rect 237 14 266 198
rect 312 14 341 198
rect 237 0 341 14
rect 397 198 502 211
rect 397 14 426 198
rect 472 14 502 198
rect 397 0 502 14
rect 558 198 662 211
rect 558 14 587 198
rect 633 14 662 198
rect 558 0 662 14
rect 718 198 806 211
rect 718 14 747 198
rect 793 14 806 198
rect 718 0 806 14
<< pdiffc >>
rect -215 14 -169 198
rect -55 14 -9 198
rect 105 14 151 198
rect 266 14 312 198
rect 426 14 472 198
rect 587 14 633 198
rect 747 14 793 198
<< polysilicon >>
rect -140 211 -84 255
rect 20 211 76 255
rect 181 211 237 255
rect 341 211 397 255
rect 502 211 558 255
rect 662 211 718 255
rect -140 -45 -84 0
rect 20 -45 76 0
rect 181 -45 237 0
rect 341 -45 397 0
rect 502 -45 558 0
rect 662 -45 718 0
<< metal1 >>
rect -215 198 -169 211
rect -215 0 -169 14
rect -55 198 -9 211
rect -55 0 -9 14
rect 105 198 151 211
rect 105 0 151 14
rect 266 198 312 211
rect 266 0 312 14
rect 426 198 472 211
rect 426 0 472 14
rect 587 198 633 211
rect 587 0 633 14
rect 747 198 793 211
rect 747 0 793 14
<< labels >>
flabel pdiffc 289 105 289 105 0 FreeSans 186 0 0 0 D
flabel pdiffc 140 105 140 105 0 FreeSans 186 0 0 0 S
flabel pdiffc -20 105 -20 105 0 FreeSans 186 0 0 0 D
flabel pdiffc -180 105 -180 105 0 FreeSans 186 0 0 0 S
flabel pdiffc 437 105 437 105 0 FreeSans 186 0 0 0 S
flabel pdiffc 598 105 598 105 0 FreeSans 186 0 0 0 D
flabel pdiffc 757 105 757 105 0 FreeSans 186 0 0 0 S
<< end >>
