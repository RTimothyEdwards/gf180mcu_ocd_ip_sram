magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal1 >>
rect -44 330 44 351
rect -44 -330 -26 330
rect 26 -330 44 330
rect -44 -351 44 -330
<< via1 >>
rect -26 -330 26 330
<< metal2 >>
rect -44 330 44 351
rect -44 -330 -26 330
rect 26 -330 44 330
rect -44 -351 44 -330
<< end >>
