magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< error_p >>
rect -75 0 -29 112
rect 85 0 131 112
<< nwell >>
rect -174 -86 230 198
<< pmos >>
rect 0 0 56 112
<< pdiff >>
rect -88 99 0 112
rect -88 13 -75 99
rect -29 13 0 99
rect -88 0 0 13
rect 56 99 144 112
rect 56 13 85 99
rect 131 13 144 99
rect 56 0 144 13
<< pdiffc >>
rect -75 13 -29 99
rect 85 13 131 99
<< polysilicon >>
rect 0 112 56 156
rect 0 -44 56 0
<< metal1 >>
rect -75 99 -29 112
rect -75 0 -29 13
rect 85 99 131 112
rect 85 0 131 13
<< labels >>
flabel pdiffc -40 56 -40 56 0 FreeSans 186 0 0 0 S
flabel pdiffc 96 56 96 56 0 FreeSans 186 0 0 0 D
<< end >>
