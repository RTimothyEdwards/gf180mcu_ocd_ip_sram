magic
tech gf180mcuD
magscale 1 10
timestamp 1764700137
<< error_s >>
rect 13150 11571 13205 11572
<< nwell >>
rect 13033 11253 13150 11572
rect 194 3187 4040 5289
rect 320 1049 3826 1666
rect 1430 1048 2963 1049
rect 4914 88 5825 603
<< pmos >>
rect 5120 186 5176 399
rect 5249 186 5305 399
rect 5434 186 5490 399
rect 5562 186 5618 399
<< pdiff >>
rect 5009 386 5120 399
rect 5009 212 5033 386
rect 5079 212 5120 386
rect 5009 186 5120 212
rect 5176 186 5249 399
rect 5305 386 5434 399
rect 5305 212 5346 386
rect 5392 212 5434 386
rect 5305 186 5434 212
rect 5490 186 5562 399
rect 5618 386 5729 399
rect 5618 212 5660 386
rect 5706 212 5729 386
rect 5618 186 5729 212
<< pdiffc >>
rect 5033 212 5079 386
rect 5346 212 5392 386
rect 5660 212 5706 386
<< psubdiff >>
rect 333 6383 12848 6418
rect 333 6337 610 6383
rect 12831 6337 12848 6383
rect 333 6302 12848 6337
<< nsubdiff >>
rect 12987 11356 13033 11469
<< psubdiffcont >>
rect 610 6337 12831 6383
<< polysilicon >>
rect 4466 531 4522 676
rect 5249 659 5289 861
rect 5433 659 5489 679
rect 5021 564 5176 623
rect 5081 558 5176 564
rect 4446 530 4522 531
rect 4383 478 4599 530
rect 4383 395 4439 478
rect 4543 395 4599 478
rect 5120 399 5176 558
rect 5249 613 5489 659
rect 5593 655 5649 657
rect 5562 640 5649 655
rect 5249 574 5490 613
rect 5249 399 5305 574
rect 5434 399 5490 574
rect 5562 569 5627 640
rect 5562 399 5618 569
rect 4383 84 4439 164
rect 4543 84 4599 164
rect 5120 135 5176 186
rect 5249 135 5305 186
rect 5434 135 5490 186
rect 5562 135 5618 186
<< metal1 >>
rect 274 11285 13029 11454
rect 279 6511 360 6512
rect 749 6511 830 6512
rect 1063 6511 1144 6512
rect 1533 6511 1614 6512
rect 1847 6511 1928 6512
rect 2317 6511 2398 6512
rect 2631 6511 2712 6512
rect 3101 6511 3182 6512
rect 3415 6511 3496 6512
rect 3885 6511 3966 6512
rect 4199 6511 4280 6512
rect 4669 6511 4750 6512
rect 4983 6511 5064 6512
rect 5453 6511 5534 6512
rect 5767 6511 5848 6512
rect 6237 6511 6318 6512
rect 6551 6511 6632 6512
rect 7021 6511 7102 6512
rect 7335 6511 7416 6512
rect 7805 6511 7886 6512
rect 8119 6511 8200 6512
rect 8589 6511 8670 6512
rect 8903 6511 8984 6512
rect 9373 6511 9454 6512
rect 9687 6511 9768 6512
rect 10157 6511 10238 6512
rect 10471 6511 10552 6512
rect 10941 6511 11022 6512
rect 11254 6511 11336 6512
rect 11725 6511 11806 6512
rect 12038 6511 12120 6512
rect 12509 6511 12590 6512
rect 12822 6511 12903 6512
rect 261 6383 12903 6511
rect 261 6337 610 6383
rect 12831 6337 12903 6383
rect 261 6087 12903 6337
rect 869 3155 959 3537
rect 3779 137 3869 1482
rect 4369 1132 4450 1183
rect 4370 949 4450 1132
rect 4369 754 4450 949
rect 4536 611 4617 826
rect 5352 707 5403 1202
rect 5517 640 5564 883
rect 5666 789 8612 1206
rect 5666 707 5721 789
rect 3933 518 4617 611
rect 5341 556 5564 640
rect 4095 196 4351 436
rect 4467 264 4516 518
rect 4633 386 5096 436
rect 4633 212 5033 386
rect 5079 212 5096 386
rect 4633 196 5096 212
rect 5015 193 5096 196
rect 5341 386 5397 556
rect 5341 212 5346 386
rect 5392 212 5397 386
rect 5341 137 5397 212
rect 5642 386 8461 476
rect 5642 212 5660 386
rect 5706 212 8461 386
rect 5642 193 8461 212
rect 3779 53 5397 137
<< metal2 >>
rect 1853 7705 1943 7989
rect 2637 7559 2727 7989
rect 3421 7492 3511 7989
rect 3420 7413 3511 7492
rect 4205 7346 4295 7989
rect 4204 7267 4295 7346
rect 4989 7200 5079 7989
rect 4407 6108 4498 7039
rect 4718 6108 4809 7200
rect 4988 7107 5079 7200
rect 5551 6108 5642 7332
rect 5773 6975 5863 7989
rect 6143 6748 6234 7479
rect 5862 6654 6234 6748
rect 5862 6108 5952 6654
rect 6695 6108 6785 7624
rect 7015 6661 7105 7770
rect 7006 6567 7105 6661
rect 7340 6678 7431 7916
rect 7800 6933 7891 8076
rect 8124 7705 8215 7989
rect 8908 7559 8999 7989
rect 9692 7413 9783 7989
rect 10476 7267 10567 7989
rect 11260 7121 11351 7989
rect 12044 6975 12135 8141
rect 7800 6840 8240 6933
rect 7340 6584 7929 6678
rect 7006 6108 7096 6567
rect 7839 6108 7929 6584
rect 8150 6108 8240 6840
rect 1229 2732 1319 3537
rect 2053 3014 2143 3537
rect 2412 2590 2503 3537
rect 3236 2873 3327 3537
rect 3596 2449 3686 3376
rect 3780 1849 4023 1943
rect 1267 424 1358 518
rect 2451 424 2541 518
rect 3635 424 3725 518
rect 3933 389 4023 1849
rect 5181 891 5271 984
rect 5002 578 5826 632
rect 5135 572 5632 578
<< metal3 >>
rect 125 9961 6479 10122
rect 12348 9961 18674 10122
rect 125 9723 5697 9884
rect 11564 9723 18674 9884
rect 125 9485 4911 9646
rect 10780 9485 18674 9646
rect 125 9247 4127 9408
rect 9996 9247 18674 9408
rect 125 9009 3343 9170
rect 9212 9009 18674 9170
rect 125 8771 2559 8932
rect 8428 8771 18674 8932
rect 125 8533 1775 8694
rect 7642 8533 18674 8694
rect 125 8295 991 8456
rect 6860 8295 18674 8456
rect 286 7997 7891 8061
rect 1069 7851 7431 7916
rect 1853 7705 8215 7770
rect 2637 7559 8999 7624
rect 3420 7413 9783 7478
rect 4204 7267 10567 7332
rect 4841 7121 11351 7186
rect 4334 6975 12135 7039
rect 268 5582 8712 6464
rect 293 1660 4108 2137
rect 310 1214 3829 1576
rect 3868 1033 4036 1137
rect 4144 1033 8612 1213
rect 3868 685 8612 1033
rect 4036 634 8612 685
rect 4144 454 8609 469
rect 3985 158 8609 454
use M1_NWELL12_3v256x8m81  M1_NWELL12_3v256x8m81_0
timestamp 1763766357
transform 1 0 6640 0 1 11412
box -6463 -159 6463 159
use M1_NWELL13_3v256x8m81  M1_NWELL13_3v256x8m81_0
timestamp 1763766357
transform 1 0 7147 0 1 309
box -1427 -216 1427 216
use M1_POLY24310591302019_3v256x8m81  M1_POLY24310591302019_3v256x8m81_0
timestamp 1764700137
transform 0 -1 5705 1 0 605
box -36 -80 36 78
use M1_POLY24310591302019_3v256x8m81  M1_POLY24310591302019_3v256x8m81_1
timestamp 1764700137
transform 1 0 5229 0 1 798
box -36 -80 36 78
use M1_POLY24310591302030_3v256x8m81  M1_POLY24310591302030_3v256x8m81_0
timestamp 1764700137
transform 1 0 4496 0 1 120
box -95 -36 95 36
use M1_POLY24310591302031_3v256x8m81  M1_POLY24310591302031_3v256x8m81_0
timestamp 1764700137
transform 1 0 5051 0 1 594
box -36 -36 36 36
use M1_PSUB$$47114284_3v256x8m81  M1_PSUB$$47114284_3v256x8m81_0
timestamp 1763766357
transform 1 0 7168 0 1 898
box -1328 -114 1328 114
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_0
timestamp 1763766357
transform -1 0 5226 0 1 861
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_1
timestamp 1763766357
transform -1 0 3978 0 1 512
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_2
timestamp 1763766357
transform -1 0 4412 0 1 826
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_3
timestamp 1763766357
transform -1 0 4857 0 1 338
box -43 -122 43 122
use M2_M1$$43375660_3v256x8m81  M2_M1$$43375660_3v256x8m81_4
timestamp 1763766357
transform -1 0 4138 0 1 325
box -43 -122 43 122
use M2_M1$$46894124_3v256x8m81  M2_M1$$46894124_3v256x8m81_0
timestamp 1764700137
transform -1 0 3641 0 1 2482
box -44 -46 45 46
use M2_M1$$46894124_3v256x8m81  M2_M1$$46894124_3v256x8m81_1
timestamp 1764700137
transform -1 0 3281 0 1 2905
box -44 -46 45 46
use M2_M1$$46894124_3v256x8m81  M2_M1$$46894124_3v256x8m81_2
timestamp 1764700137
transform -1 0 1274 0 1 2764
box -44 -46 45 46
use M2_M1$$46894124_3v256x8m81  M2_M1$$46894124_3v256x8m81_3
timestamp 1764700137
transform -1 0 2457 0 1 2622
box -44 -46 45 46
use M2_M1$$46894124_3v256x8m81  M2_M1$$46894124_3v256x8m81_4
timestamp 1764700137
transform -1 0 2098 0 1 3047
box -44 -46 45 46
use M2_M1$$47630380_3v256x8m81  M2_M1$$47630380_3v256x8m81_0
timestamp 1763766357
transform -1 0 7016 0 1 334
box -1373 -123 1373 123
use M2_M1$$47631404_3v256x8m81  M2_M1$$47631404_3v256x8m81_0
timestamp 1763766357
transform -1 0 7109 0 1 919
box -1299 -123 1299 123
use M2_M14310591302051_3v256x8m81  M2_M14310591302051_3v256x8m81_0
timestamp 1763766357
transform 1 0 5047 0 1 605
box -99 -34 99 34
use M2_M14310591302051_3v256x8m81  M2_M14310591302051_3v256x8m81_1
timestamp 1763766357
transform 1 0 5727 0 1 605
box -99 -34 99 34
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_0
timestamp 1763766357
transform -1 0 4412 0 1 826
box -44 -123 44 123
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_1
timestamp 1763766357
transform -1 0 4857 0 1 338
box -44 -123 44 123
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_2
timestamp 1763766357
transform -1 0 4138 0 1 325
box -44 -123 44 123
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_3
timestamp 1763766357
transform 1 0 1898 0 1 7647
box -44 -123 44 123
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_4
timestamp 1763766357
transform 1 0 330 0 1 8018
box -44 -123 44 123
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_5
timestamp 1763766357
transform 1 0 7845 0 1 8029
box -44 -123 44 123
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_6
timestamp 1763766357
transform 1 0 8954 0 1 7682
box -44 -123 44 123
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_7
timestamp 1763766357
transform 1 0 9738 0 1 7536
box -44 -123 44 123
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_8
timestamp 1763766357
transform 1 0 10522 0 1 7389
box -44 -123 44 123
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_9
timestamp 1763766357
transform 1 0 11306 0 1 7244
box -44 -123 44 123
use M3_M2$$43368492_3v256x8m81  M3_M2$$43368492_3v256x8m81_10
timestamp 1763766357
transform 1 0 12090 0 1 7098
box -44 -123 44 123
use M3_M2$$43368492_R90_3v256x8m81  M3_M2$$43368492_R90_3v256x8m81_0
timestamp 1764700137
transform 0 -1 7459 1 0 7883
box -46 -119 46 119
use M3_M2$$43368492_R270_3v256x8m81  M3_M2$$43368492_R270_3v256x8m81_0
timestamp 1763766357
transform 0 1 8243 -1 0 7742
box -46 -119 46 119
use M3_M2$$43371564_3v256x8m81  M3_M2$$43371564_3v256x8m81_0
timestamp 1764700137
transform 1 0 6188 0 1 7445
box -119 -46 119 46
use M3_M2$$43371564_3v256x8m81  M3_M2$$43371564_3v256x8m81_1
timestamp 1764700137
transform 1 0 4899 0 1 7154
box -119 -46 119 46
use M3_M2$$43371564_3v256x8m81  M3_M2$$43371564_3v256x8m81_2
timestamp 1764700137
transform 1 0 4453 0 1 7007
box -119 -46 119 46
use M3_M2$$43371564_3v256x8m81  M3_M2$$43371564_3v256x8m81_3
timestamp 1764700137
transform 1 0 5891 0 1 7007
box -119 -46 119 46
use M3_M2$$43371564_3v256x8m81  M3_M2$$43371564_3v256x8m81_4
timestamp 1764700137
transform 1 0 5523 0 1 7299
box -119 -46 119 46
use M3_M2$$43371564_3v256x8m81  M3_M2$$43371564_3v256x8m81_5
timestamp 1764700137
transform 1 0 4250 0 1 7299
box -119 -46 119 46
use M3_M2$$43371564_3v256x8m81  M3_M2$$43371564_3v256x8m81_6
timestamp 1764700137
transform 1 0 3466 0 1 7445
box -119 -46 119 46
use M3_M2$$43371564_3v256x8m81  M3_M2$$43371564_3v256x8m81_7
timestamp 1764700137
transform 1 0 2755 0 1 7591
box -119 -46 119 46
use M3_M2$$43371564_3v256x8m81  M3_M2$$43371564_3v256x8m81_8
timestamp 1764700137
transform 1 0 1188 0 1 7883
box -119 -46 119 46
use M3_M2$$43371564_3v256x8m81  M3_M2$$43371564_3v256x8m81_9
timestamp 1764700137
transform 1 0 6666 0 1 7591
box -119 -46 119 46
use M3_M2$$43371564_3v256x8m81  M3_M2$$43371564_3v256x8m81_10
timestamp 1764700137
transform 1 0 6675 0 1 8062
box -119 -46 119 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_0
timestamp 1764700137
transform 1 0 6434 0 1 10042
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_1
timestamp 1764700137
transform 1 0 6120 0 1 10042
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_2
timestamp 1764700137
transform 1 0 633 0 1 8375
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_3
timestamp 1764700137
transform 1 0 947 0 1 8375
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_4
timestamp 1764700137
transform 1 0 1731 0 1 8613
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_5
timestamp 1764700137
transform 1 0 1417 0 1 8613
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_6
timestamp 1764700137
transform 1 0 2515 0 1 8851
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_7
timestamp 1764700137
transform 1 0 2201 0 1 8851
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_8
timestamp 1764700137
transform 1 0 3299 0 1 9089
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_9
timestamp 1764700137
transform 1 0 2985 0 1 9089
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_10
timestamp 1764700137
transform 1 0 4083 0 1 9327
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_11
timestamp 1764700137
transform 1 0 3769 0 1 9327
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_12
timestamp 1764700137
transform 1 0 4867 0 1 9565
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_13
timestamp 1764700137
transform 1 0 4553 0 1 9565
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_14
timestamp 1764700137
transform 1 0 5650 0 1 9804
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_15
timestamp 1764700137
transform 1 0 5337 0 1 9804
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_16
timestamp 1764700137
transform -1 0 7218 0 -1 8375
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_17
timestamp 1764700137
transform -1 0 6904 0 -1 8375
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_18
timestamp 1764700137
transform -1 0 8002 0 -1 8613
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_19
timestamp 1764700137
transform -1 0 7688 0 -1 8613
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_20
timestamp 1764700137
transform -1 0 8786 0 -1 8851
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_21
timestamp 1764700137
transform -1 0 8472 0 -1 8851
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_22
timestamp 1764700137
transform -1 0 9570 0 -1 9089
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_23
timestamp 1764700137
transform -1 0 9256 0 -1 9089
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_24
timestamp 1764700137
transform -1 0 10354 0 -1 9327
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_25
timestamp 1764700137
transform -1 0 10040 0 -1 9327
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_26
timestamp 1764700137
transform -1 0 11138 0 -1 9565
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_27
timestamp 1764700137
transform -1 0 10824 0 -1 9565
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_28
timestamp 1764700137
transform -1 0 11922 0 -1 9804
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_29
timestamp 1764700137
transform -1 0 11608 0 -1 9804
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_30
timestamp 1764700137
transform -1 0 12392 0 -1 10042
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_31
timestamp 1764700137
transform -1 0 12706 0 -1 10042
box -45 -46 45 46
use M3_M2$$46895148_3v256x8m81  M3_M2$$46895148_3v256x8m81_32
timestamp 1764700137
transform 1 0 7060 0 1 7737
box -45 -46 45 46
use M3_M2$$47632428_3v256x8m81  M3_M2$$47632428_3v256x8m81_0
timestamp 1763766357
transform -1 0 7016 0 1 334
box -1373 -123 1373 123
use M3_M2$$47633452_3v256x8m81  M3_M2$$47633452_3v256x8m81_0
timestamp 1763766357
transform -1 0 7109 0 1 919
box -1299 -123 1299 123
use nmos_1p2$$47342636_3v256x8m81  nmos_1p2$$47342636_3v256x8m81_0
timestamp 1763766357
transform -1 0 4508 0 1 697
box -102 -44 130 170
use nmos_5p04310591302056_3v256x8m81  nmos_5p04310591302056_3v256x8m81_0
timestamp 1763766357
transform -1 0 5489 0 1 701
box -88 -44 144 222
use nmos_5p04310591302056_3v256x8m81  nmos_5p04310591302056_3v256x8m81_1
timestamp 1763766357
transform -1 0 5649 0 1 701
box -88 -44 144 222
use pmos_1p2$$47109164_3v256x8m81  pmos_1p2$$47109164_3v256x8m81_0
timestamp 1763766357
transform -1 0 4557 0 1 196
box -216 -86 348 245
use ypredec1_bot_3v256x8m81  ypredec1_bot_3v256x8m81_0
timestamp 1764700137
transform 1 0 2636 0 1 718
box -14 -33 1367 5518
use ypredec1_bot_3v256x8m81  ypredec1_bot_3v256x8m81_1
timestamp 1764700137
transform 1 0 268 0 1 718
box -14 -33 1367 5518
use ypredec1_bot_3v256x8m81  ypredec1_bot_3v256x8m81_2
timestamp 1764700137
transform 1 0 1452 0 1 718
box -14 -33 1367 5518
use ypredec1_xax8_3v256x8m81  ypredec1_xax8_3v256x8m81_0
timestamp 1764700137
transform 1 0 3936 0 1 1069
box -1 -38 4792 5176
use ypredec1_ys_3v256x8m81  ypredec1_ys_3v256x8m81_0
timestamp 1764700137
transform 1 0 2530 0 1 6337
box 0 0 1351 5167
use ypredec1_ys_3v256x8m81  ypredec1_ys_3v256x8m81_1
timestamp 1764700137
transform 1 0 3314 0 1 6337
box 0 0 1351 5167
use ypredec1_ys_3v256x8m81  ypredec1_ys_3v256x8m81_2
timestamp 1764700137
transform 1 0 4098 0 1 6337
box 0 0 1351 5167
use ypredec1_ys_3v256x8m81  ypredec1_ys_3v256x8m81_3
timestamp 1764700137
transform 1 0 4882 0 1 6337
box 0 0 1351 5167
use ypredec1_ys_3v256x8m81  ypredec1_ys_3v256x8m81_4
timestamp 1764700137
transform 1 0 178 0 1 6337
box 0 0 1351 5167
use ypredec1_ys_3v256x8m81  ypredec1_ys_3v256x8m81_5
timestamp 1764700137
transform 1 0 962 0 1 6337
box 0 0 1351 5167
use ypredec1_ys_3v256x8m81  ypredec1_ys_3v256x8m81_6
timestamp 1764700137
transform 1 0 1746 0 1 6337
box 0 0 1351 5167
use ypredec1_ys_3v256x8m81  ypredec1_ys_3v256x8m81_7
timestamp 1764700137
transform 1 0 10370 0 1 6337
box 0 0 1351 5167
use ypredec1_ys_3v256x8m81  ypredec1_ys_3v256x8m81_8
timestamp 1764700137
transform 1 0 11154 0 1 6337
box 0 0 1351 5167
use ypredec1_ys_3v256x8m81  ypredec1_ys_3v256x8m81_9
timestamp 1764700137
transform 1 0 11938 0 1 6337
box 0 0 1351 5167
use ypredec1_ys_3v256x8m81  ypredec1_ys_3v256x8m81_10
timestamp 1764700137
transform 1 0 7234 0 1 6337
box 0 0 1351 5167
use ypredec1_ys_3v256x8m81  ypredec1_ys_3v256x8m81_11
timestamp 1764700137
transform 1 0 8018 0 1 6337
box 0 0 1351 5167
use ypredec1_ys_3v256x8m81  ypredec1_ys_3v256x8m81_12
timestamp 1764700137
transform 1 0 8802 0 1 6337
box 0 0 1351 5167
use ypredec1_ys_3v256x8m81  ypredec1_ys_3v256x8m81_13
timestamp 1764700137
transform 1 0 9586 0 1 6337
box 0 0 1351 5167
use ypredec1_ys_3v256x8m81  ypredec1_ys_3v256x8m81_14
timestamp 1764700137
transform 1 0 6450 0 1 6337
box 0 0 1351 5167
use ypredec1_ys_3v256x8m81  ypredec1_ys_3v256x8m81_15
timestamp 1764700137
transform 1 0 5666 0 1 6337
box 0 0 1351 5167
<< labels >>
rlabel metal3 s 695 9565 695 9565 4 ly[5]
port 1 nsew
rlabel metal3 s 695 9327 695 9327 4 ly[4]
port 2 nsew
rlabel metal3 s 695 10042 695 10042 4 ly[7]
port 3 nsew
rlabel metal3 s 695 9089 695 9089 4 ly[3]
port 4 nsew
rlabel metal3 s 695 8851 695 8851 4 ly[2]
port 5 nsew
rlabel metal3 s 695 8613 695 8613 4 ly[1]
port 6 nsew
rlabel metal3 s 695 8375 695 8375 4 ly[0]
port 7 nsew
rlabel metal3 s 17875 8375 17875 8375 4 ry[0]
port 8 nsew
rlabel metal3 s 17875 8613 17875 8613 4 ry[1]
port 9 nsew
rlabel metal3 s 17875 8851 17875 8851 4 ry[2]
port 10 nsew
rlabel metal3 s 17875 9089 17875 9089 4 ry[3]
port 11 nsew
rlabel metal3 s 17875 9327 17875 9327 4 ry[4]
port 12 nsew
rlabel metal3 s 17875 9565 17875 9565 4 ry[5]
port 13 nsew
rlabel metal3 s 17875 9804 17875 9804 4 ry[6]
port 14 nsew
rlabel metal3 s 17875 10042 17875 10042 4 ry[7]
port 15 nsew
rlabel metal3 s 695 9804 695 9804 4 ly[6]
port 16 nsew
rlabel metal2 s 5819 598 5819 598 4 men
port 17 nsew
rlabel metal2 s 3679 471 3679 471 4 A[0]
port 18 nsew
rlabel metal2 s 2496 471 2496 471 4 A[1]
port 19 nsew
rlabel metal2 s 1312 471 1312 471 4 A[2]
port 20 nsew
rlabel metal2 s 5226 934 5226 934 4 clk
port 21 nsew
<< end >>
