magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal2 >>
rect -113 323 113 330
rect -113 -323 -106 323
rect 106 -323 113 323
rect -113 -330 113 -323
<< via2 >>
rect -106 -323 106 323
<< metal3 >>
rect -113 323 113 330
rect -113 -323 -106 323
rect 106 -323 113 323
rect -113 -330 113 -323
<< end >>
