magic
tech gf180mcuD
magscale 1 10
timestamp 1764623439
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_0
timestamp 1764525316
transform 1 0 3194 0 1 1978
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_1
timestamp 1764525316
transform 1 0 2723 0 1 1978
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_2
timestamp 1764525316
transform 1 0 280 0 1 2118
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_3
timestamp 1764525316
transform 1 0 1064 0 1 2118
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_4
timestamp 1764525316
transform 1 0 4024 0 1 1836
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_5
timestamp 1764525316
transform 1 0 4181 0 1 1412
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_6
timestamp 1764525316
transform 1 0 750 0 1 1412
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_7
timestamp 1764525316
transform 1 0 593 0 1 1836
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_8
timestamp 1764525316
transform 1 0 3350 0 1 1694
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_9
timestamp 1764525316
transform 1 0 2566 0 1 1694
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_10
timestamp 1764525316
transform 1 0 3867 0 1 1553
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_11
timestamp 1764525316
transform 1 0 4337 0 1 1553
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_12
timestamp 1764525316
transform 1 0 2050 0 1 1553
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_13
timestamp 1764525316
transform 1 0 1579 0 1 1553
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_14
timestamp 1764525316
transform 1 0 1893 0 1 1412
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_15
timestamp 1764525316
transform 1 0 1736 0 1 1836
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_16
timestamp 1764525316
transform 1 0 4494 0 1 1694
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_17
timestamp 1764525316
transform 1 0 2207 0 1 2118
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_18
timestamp 1764525316
transform 1 0 1423 0 1 2118
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_19
timestamp 1764525316
transform 1 0 3710 0 1 1694
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_20
timestamp 1764525316
transform 1 0 907 0 1 1978
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_21
timestamp 1764525316
transform 1 0 436 0 1 1978
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_22
timestamp 1764525316
transform 1 0 2880 0 1 1836
box -67 -48 67 47
use M1_POLY2$$44753964_3v512x8m81  M1_POLY2$$44753964_3v512x8m81_23
timestamp 1764525316
transform 1 0 3037 0 1 1412
box -67 -48 67 47
use M2_M14310591302057_3v512x8m81  M2_M14310591302057_3v512x8m81_0
timestamp 1764525316
transform 1 0 1815 0 1 701
box -34 -354 34 354
use M2_M14310591302057_3v512x8m81  M2_M14310591302057_3v512x8m81_1
timestamp 1764525316
transform 1 0 2958 0 1 701
box -34 -354 34 354
use M2_M14310591302057_3v512x8m81  M2_M14310591302057_3v512x8m81_2
timestamp 1764525316
transform 1 0 4102 0 1 701
box -34 -354 34 354
use M2_M14310591302057_3v512x8m81  M2_M14310591302057_3v512x8m81_3
timestamp 1764525316
transform 1 0 672 0 1 701
box -34 -354 34 354
use M3_M24310591302058_3v512x8m81  M3_M24310591302058_3v512x8m81_0
timestamp 1764525316
transform 1 0 672 0 1 701
box -35 -354 35 354
use M3_M24310591302058_3v512x8m81  M3_M24310591302058_3v512x8m81_1
timestamp 1764525316
transform 1 0 2958 0 1 701
box -35 -354 35 354
use M3_M24310591302058_3v512x8m81  M3_M24310591302058_3v512x8m81_2
timestamp 1764525316
transform 1 0 4102 0 1 701
box -35 -354 35 354
use M3_M24310591302058_3v512x8m81  M3_M24310591302058_3v512x8m81_3
timestamp 1764525316
transform 1 0 1815 0 1 701
box -35 -354 35 354
use ypredec1_xa_3v512x8m81  ypredec1_xa_3v512x8m81_0
timestamp 1764525316
transform -1 0 3060 0 1 4948
box -100 -4986 774 228
use ypredec1_xa_3v512x8m81  ypredec1_xa_3v512x8m81_1
timestamp 1764525316
transform -1 0 4204 0 1 4948
box -100 -4986 774 228
use ypredec1_xa_3v512x8m81  ypredec1_xa_3v512x8m81_2
timestamp 1764525316
transform -1 0 1916 0 1 4948
box -100 -4986 774 228
use ypredec1_xa_3v512x8m81  ypredec1_xa_3v512x8m81_3
timestamp 1764525316
transform -1 0 773 0 1 4948
box -100 -4986 774 228
use ypredec1_xa_3v512x8m81  ypredec1_xa_3v512x8m81_4
timestamp 1764525316
transform 1 0 2874 0 1 4948
box -100 -4986 774 228
use ypredec1_xa_3v512x8m81  ypredec1_xa_3v512x8m81_5
timestamp 1764525316
transform 1 0 4018 0 1 4948
box -100 -4986 774 228
use ypredec1_xa_3v512x8m81  ypredec1_xa_3v512x8m81_6
timestamp 1764525316
transform 1 0 1730 0 1 4948
box -100 -4986 774 228
use ypredec1_xa_3v512x8m81  ypredec1_xa_3v512x8m81_7
timestamp 1764525316
transform 1 0 587 0 1 4948
box -100 -4986 774 228
<< properties >>
string MASKHINTS_PPLUS 132 2192 4659 2813 132 3755 4659 4385
<< end >>
