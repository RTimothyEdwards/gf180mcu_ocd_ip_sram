magic
tech gf180mcuD
magscale 1 10
timestamp 1765925964
<< metal1 >>
rect 401 77537 447 77650
rect 401 76769 447 76882
rect 401 76325 447 76438
rect 401 75557 447 75670
rect 401 75113 447 75226
rect 401 74345 447 74458
rect 401 73901 447 74014
rect 401 73133 447 73246
rect 401 72689 447 72802
rect 401 71921 447 72034
rect 401 71477 447 71590
rect 401 70709 447 70822
rect 401 70265 447 70378
rect 401 69497 447 69610
rect 401 69053 447 69166
rect 401 68285 447 68398
rect 401 67841 447 67954
rect 401 67073 447 67186
rect 401 66629 447 66742
rect 401 65861 447 65974
rect 401 65417 447 65530
rect 401 64649 447 64762
rect 401 64205 447 64318
rect 401 63437 447 63550
rect 401 62993 447 63106
rect 401 62225 447 62338
rect 401 61781 447 61894
rect 401 61013 447 61126
rect 401 60569 447 60682
rect 401 59801 447 59914
rect 401 59357 447 59470
rect 401 58589 447 58702
rect 401 58145 447 58258
rect 401 57377 447 57490
rect 401 56933 447 57046
rect 401 56165 447 56278
rect 401 55721 447 55834
rect 401 54953 447 55066
rect 401 54509 447 54622
rect 401 53741 447 53854
rect 401 53297 447 53410
rect 401 52529 447 52642
rect 401 52085 447 52198
rect 401 51317 447 51430
rect 401 50873 447 50986
rect 401 50105 447 50218
rect 401 49661 447 49774
rect 401 48893 447 49006
rect 401 48449 447 48562
rect 401 47681 447 47794
rect 401 47237 447 47350
rect 401 46469 447 46582
rect 401 46025 447 46138
rect 401 45257 447 45370
rect 401 44813 447 44926
rect 401 44045 447 44158
rect 401 43601 447 43714
rect 401 42833 447 42946
rect 401 42389 447 42502
rect 401 41621 447 41734
rect 401 41177 447 41290
rect 401 40409 447 40522
rect 401 39965 447 40078
rect 401 39197 447 39310
rect 401 38753 447 38866
rect 401 37985 447 38098
rect 401 37541 447 37654
rect 401 36773 447 36886
rect 401 36329 447 36442
rect 401 35561 447 35674
rect 401 35117 447 35230
rect 401 34349 447 34462
rect 401 33905 447 34018
rect 401 33137 447 33250
rect 401 32693 447 32806
rect 401 31925 447 32038
rect 401 31481 447 31594
rect 401 30713 447 30826
rect 401 30269 447 30382
rect 401 29501 447 29614
rect 401 29057 447 29170
rect 401 28289 447 28402
rect 401 27845 447 27958
rect 401 27077 447 27190
rect 401 26633 447 26746
rect 401 25865 447 25978
rect 401 25421 447 25534
rect 401 24653 447 24766
rect 401 24209 447 24322
rect 401 23441 447 23554
rect 401 22997 447 23110
rect 401 22229 447 22342
rect 401 21785 447 21898
rect 401 21017 447 21130
rect 401 20573 447 20686
rect 401 19805 447 19918
rect 401 19361 447 19474
rect 401 18593 447 18706
rect 401 18149 447 18262
rect 401 17381 447 17494
rect 401 16937 447 17050
rect 401 16169 447 16282
rect 401 15725 447 15838
rect 401 14957 447 15070
rect 401 14513 447 14626
rect 401 13745 447 13858
rect 401 13301 447 13414
rect 401 12533 447 12646
rect 401 12089 447 12202
rect 401 11321 447 11434
rect 401 10877 447 10990
rect 401 10109 447 10222
rect 401 9665 447 9778
rect 401 8897 447 9010
rect 401 8453 447 8566
rect 401 7685 447 7798
rect 401 7241 447 7354
rect 401 6473 447 6586
rect 401 6029 447 6142
rect 401 5261 447 5374
rect 401 4817 447 4930
rect 401 4049 447 4162
rect 401 3605 447 3718
rect 401 2837 447 2950
rect 401 2393 447 2506
rect 401 1625 447 1738
rect 401 1181 447 1294
rect 401 413 447 526
<< metal2 >>
rect 734 129 854 229
rect 946 129 1066 229
rect 1170 129 1290 229
rect 1382 129 1502 229
rect 1606 129 1726 229
rect 1818 129 1938 229
rect 2042 129 2162 229
rect 2254 129 2374 229
rect 2478 129 2598 229
rect 2690 129 2810 229
rect 2914 129 3034 229
rect 3126 129 3246 229
rect 3350 129 3470 229
rect 3562 129 3682 229
rect 3786 129 3906 229
rect 3998 129 4118 229
rect 4642 129 4762 229
rect 4854 129 4974 229
rect 5078 129 5198 229
rect 5290 129 5410 229
rect 5514 129 5634 229
rect 5726 129 5846 229
rect 5950 129 6070 229
rect 6162 129 6282 229
rect 6386 129 6506 229
rect 6598 129 6718 229
rect 6822 129 6942 229
rect 7034 129 7154 229
rect 7258 129 7378 229
rect 7470 129 7590 229
rect 7694 129 7814 229
rect 7906 129 8026 229
rect 8550 129 8670 229
rect 8762 129 8882 229
rect 8986 129 9106 229
rect 9198 129 9318 229
rect 9422 129 9542 229
rect 9634 129 9754 229
rect 9858 129 9978 229
rect 10070 129 10190 229
rect 10294 129 10414 229
rect 10506 129 10626 229
rect 10730 129 10850 229
rect 10942 129 11062 229
rect 11166 129 11286 229
rect 11378 129 11498 229
rect 11602 129 11722 229
rect 11814 129 11934 229
rect 12458 129 12578 229
rect 12670 129 12790 229
rect 12894 129 13014 229
rect 13106 129 13226 229
rect 13330 129 13450 229
rect 13542 129 13662 229
rect 13766 129 13886 229
rect 13978 129 14098 229
rect 14202 129 14322 229
rect 14414 129 14534 229
rect 14638 129 14758 229
rect 14850 129 14970 229
rect 15074 129 15194 229
rect 15286 129 15406 229
rect 15510 129 15630 229
rect 15722 129 15842 229
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_0
array 0 7 -436 0 63 1212
timestamp 1764626446
transform -1 0 12924 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_1
array 0 7 -436 0 63 1212
timestamp 1764626446
transform -1 0 5108 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_2
array 0 7 436 0 63 1212
timestamp 1764626446
transform 1 0 600 0 1 0
box 30 103 570 1445
use 018SRAM_cell1_2x_3v1024x8m81  018SRAM_cell1_2x_3v1024x8m81_3
array 0 7 436 0 63 1212
timestamp 1764626446
transform 1 0 8416 0 1 0
box 30 103 570 1445
use 018SRAM_strap1_2x_3v1024x8m81  018SRAM_strap1_2x_3v1024x8m81_0
array 0 0 -420 0 63 1212
timestamp 1764693440
transform -1 0 12497 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_2x_3v1024x8m81  018SRAM_strap1_2x_3v1024x8m81_1
array 0 0 -420 0 63 1212
timestamp 1764693440
transform -1 0 773 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_2x_3v1024x8m81  018SRAM_strap1_2x_3v1024x8m81_2
array 0 0 -420 0 63 1212
timestamp 1764693440
transform -1 0 4681 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_2x_3v1024x8m81  018SRAM_strap1_2x_3v1024x8m81_3
array 0 0 -420 0 63 1212
timestamp 1764693440
transform -1 0 8589 0 1 900
box 91 -797 511 545
use 018SRAM_strap1_2x_bndry_3v1024x8m81  018SRAM_strap1_2x_bndry_3v1024x8m81_0
array 0 0 420 0 63 1212
timestamp 1764625442
transform 1 0 15803 0 1 900
box 91 -797 511 545
<< labels >>
rlabel metal1 420 468 420 468 4 wl[0]
rlabel metal1 420 1236 420 1236 4 wl[1]
rlabel metal1 420 1680 420 1680 4 wl[2]
rlabel metal1 420 2448 420 2448 4 wl[3]
rlabel metal1 420 2892 420 2892 4 wl[4]
rlabel metal1 420 3660 420 3660 4 wl[5]
rlabel metal1 420 4104 420 4104 4 wl[6]
rlabel metal1 420 4872 420 4872 4 wl[7]
rlabel metal1 420 5316 420 5316 4 wl[8]
rlabel metal1 420 6084 420 6084 4 wl[9]
rlabel metal1 420 6528 420 6528 4 wl[10]
rlabel metal1 420 7296 420 7296 4 wl[11]
rlabel metal1 420 7740 420 7740 4 wl[12]
rlabel metal1 420 8508 420 8508 4 wl[13]
rlabel metal1 420 8952 420 8952 4 wl[14]
rlabel metal1 420 9720 420 9720 4 wl[15]
rlabel metal1 420 10164 420 10164 4 wl[16]
rlabel metal1 420 10932 420 10932 4 wl[17]
rlabel metal1 420 11376 420 11376 4 wl[18]
rlabel metal1 420 12144 420 12144 4 wl[19]
rlabel metal1 420 12588 420 12588 4 wl[20]
rlabel metal1 420 13356 420 13356 4 wl[21]
rlabel metal1 420 13800 420 13800 4 wl[22]
rlabel metal1 420 14568 420 14568 4 wl[23]
rlabel metal1 420 15012 420 15012 4 wl[24]
rlabel metal1 420 15780 420 15780 4 wl[25]
rlabel metal1 420 16224 420 16224 4 wl[26]
rlabel metal1 420 16992 420 16992 4 wl[27]
rlabel metal1 420 17436 420 17436 4 wl[28]
rlabel metal1 420 18204 420 18204 4 wl[29]
rlabel metal1 420 18648 420 18648 4 wl[30]
rlabel metal1 420 19416 420 19416 4 wl[31]
rlabel metal1 420 19860 420 19860 4 wl[32]
rlabel metal1 420 20628 420 20628 4 wl[33]
rlabel metal1 420 21072 420 21072 4 wl[34]
rlabel metal1 420 21840 420 21840 4 wl[35]
rlabel metal1 420 22284 420 22284 4 wl[36]
rlabel metal1 420 23052 420 23052 4 wl[37]
rlabel metal1 420 23496 420 23496 4 wl[38]
rlabel metal1 420 24264 420 24264 4 wl[39]
rlabel metal1 420 24708 420 24708 4 wl[40]
rlabel metal1 420 25476 420 25476 4 wl[41]
rlabel metal1 420 25920 420 25920 4 wl[42]
rlabel metal1 420 26688 420 26688 4 wl[43]
rlabel metal1 420 27132 420 27132 4 wl[44]
rlabel metal1 420 27900 420 27900 4 wl[45]
rlabel metal1 420 28344 420 28344 4 wl[46]
rlabel metal1 420 29112 420 29112 4 wl[47]
rlabel metal1 420 29556 420 29556 4 wl[48]
rlabel metal1 420 30324 420 30324 4 wl[49]
rlabel metal1 420 30768 420 30768 4 wl[50]
rlabel metal1 420 31536 420 31536 4 wl[51]
rlabel metal1 420 31980 420 31980 4 wl[52]
rlabel metal1 420 32748 420 32748 4 wl[53]
rlabel metal1 420 33192 420 33192 4 wl[54]
rlabel metal1 420 33960 420 33960 4 wl[55]
rlabel metal1 420 34404 420 34404 4 wl[56]
rlabel metal1 420 35172 420 35172 4 wl[57]
rlabel metal1 420 35616 420 35616 4 wl[58]
rlabel metal1 420 36384 420 36384 4 wl[59]
rlabel metal1 420 36828 420 36828 4 wl[60]
rlabel metal1 420 37596 420 37596 4 wl[61]
rlabel metal1 420 38040 420 38040 4 wl[62]
rlabel metal1 420 38808 420 38808 4 wl[63]
rlabel metal1 420 39252 420 39252 4 wl[64]
rlabel metal1 420 40020 420 40020 4 wl[65]
rlabel metal1 420 40464 420 40464 4 wl[66]
rlabel metal1 420 41232 420 41232 4 wl[67]
rlabel metal1 420 41676 420 41676 4 wl[68]
rlabel metal1 420 42444 420 42444 4 wl[69]
rlabel metal1 420 42888 420 42888 4 wl[70]
rlabel metal1 420 43656 420 43656 4 wl[71]
rlabel metal1 420 44100 420 44100 4 wl[72]
rlabel metal1 420 44868 420 44868 4 wl[73]
rlabel metal1 420 45312 420 45312 4 wl[74]
rlabel metal1 420 46080 420 46080 4 wl[75]
rlabel metal1 420 46524 420 46524 4 wl[76]
rlabel metal1 420 47292 420 47292 4 wl[77]
rlabel metal1 420 47736 420 47736 4 wl[78]
rlabel metal1 420 48504 420 48504 4 wl[79]
rlabel metal1 420 48948 420 48948 4 wl[80]
rlabel metal1 420 49716 420 49716 4 wl[81]
rlabel metal1 420 50160 420 50160 4 wl[82]
rlabel metal1 420 50928 420 50928 4 wl[83]
rlabel metal1 420 51372 420 51372 4 wl[84]
rlabel metal1 420 52140 420 52140 4 wl[85]
rlabel metal1 420 52584 420 52584 4 wl[86]
rlabel metal1 420 53352 420 53352 4 wl[87]
rlabel metal1 420 53796 420 53796 4 wl[88]
rlabel metal1 420 54564 420 54564 4 wl[89]
rlabel metal1 420 55008 420 55008 4 wl[90]
rlabel metal1 420 55776 420 55776 4 wl[91]
rlabel metal1 420 56220 420 56220 4 wl[92]
rlabel metal1 420 56988 420 56988 4 wl[93]
rlabel metal1 420 57432 420 57432 4 wl[94]
rlabel metal1 420 58200 420 58200 4 wl[95]
rlabel metal1 420 58644 420 58644 4 wl[96]
rlabel metal1 420 59412 420 59412 4 wl[97]
rlabel metal1 420 59856 420 59856 4 wl[98]
rlabel metal1 420 60624 420 60624 4 wl[99]
rlabel metal1 420 61068 420 61068 4 wl[100]
rlabel metal1 420 61836 420 61836 4 wl[101]
rlabel metal1 420 62280 420 62280 4 wl[102]
rlabel metal1 420 63048 420 63048 4 wl[103]
rlabel metal1 420 63492 420 63492 4 wl[104]
rlabel metal1 420 64260 420 64260 4 wl[105]
rlabel metal1 420 64704 420 64704 4 wl[106]
rlabel metal1 420 65472 420 65472 4 wl[107]
rlabel metal1 420 65916 420 65916 4 wl[108]
rlabel metal1 420 66684 420 66684 4 wl[109]
rlabel metal1 420 67128 420 67128 4 wl[110]
rlabel metal1 420 67896 420 67896 4 wl[111]
rlabel metal1 420 68340 420 68340 4 wl[112]
rlabel metal1 420 69108 420 69108 4 wl[113]
rlabel metal1 420 69552 420 69552 4 wl[114]
rlabel metal1 420 70320 420 70320 4 wl[115]
rlabel metal1 420 70764 420 70764 4 wl[116]
rlabel metal1 420 71532 420 71532 4 wl[117]
rlabel metal1 420 71976 420 71976 4 wl[118]
rlabel metal1 420 72744 420 72744 4 wl[119]
rlabel metal1 420 73188 420 73188 4 wl[120]
rlabel metal1 420 73956 420 73956 4 wl[121]
rlabel metal1 420 74400 420 74400 4 wl[122]
rlabel metal1 420 75168 420 75168 4 wl[123]
rlabel metal1 420 75612 420 75612 4 wl[124]
rlabel metal1 420 76380 420 76380 4 wl[125]
rlabel metal1 420 76824 420 76824 4 wl[126]
rlabel metal1 420 77592 420 77592 4 wl[127]
rlabel metal2 15349 181 15349 181 6 bb[1]
rlabel metal2 15137 181 15137 181 6 b[1]
rlabel metal2 14477 181 14477 181 6 bb[3]
rlabel metal2 14265 181 14265 181 6 b[3]
rlabel metal2 13605 181 13605 181 6 bb[5]
rlabel metal2 13393 181 13393 181 6 b[5]
rlabel metal2 12733 181 12733 181 6 bb[7]
rlabel metal2 12521 181 12521 181 6 b[7]
rlabel metal2 11437 175 11437 175 6 bb[9]
rlabel metal2 11225 175 11225 175 6 b[9]
rlabel metal2 10565 175 10565 175 6 bb[11]
rlabel metal2 10353 175 10353 175 6 b[11]
rlabel metal2 9693 175 9693 175 6 bb[13]
rlabel metal2 9481 175 9481 175 6 b[13]
rlabel metal2 8821 175 8821 175 6 bb[15]
rlabel metal2 8609 175 8609 175 6 b[15]
rlabel metal2 7531 177 7531 177 6 bb[17]
rlabel metal2 7319 177 7319 177 6 b[17]
rlabel metal2 6659 177 6659 177 6 bb[19]
rlabel metal2 6447 177 6447 177 6 b[19]
rlabel metal2 5787 177 5787 177 6 bb[21]
rlabel metal2 5575 177 5575 177 6 b[21]
rlabel metal2 4915 177 4915 177 6 bb[23]
rlabel metal2 4703 177 4703 177 6 b[23]
rlabel metal2 3623 173 3623 173 6 bb[25]
rlabel metal2 3411 173 3411 173 6 b[25]
rlabel metal2 2751 173 2751 173 6 bb[27]
rlabel metal2 2539 173 2539 173 6 b[27]
rlabel metal2 1879 173 1879 173 6 bb[29]
rlabel metal2 1667 173 1667 173 6 b[29]
rlabel metal2 1007 173 1007 173 6 bb[31]
rlabel metal2 795 173 795 173 6 b[31]
rlabel metal2 1231 173 1231 173 4 bb[30]
rlabel metal2 1443 173 1443 173 4 b[30]
rlabel metal2 2103 173 2103 173 4 bb[28]
rlabel metal2 2315 173 2315 173 4 b[28]
rlabel metal2 2975 173 2975 173 4 bb[26]
rlabel metal2 3187 173 3187 173 4 b[26]
rlabel metal2 3847 173 3847 173 4 bb[24]
rlabel metal2 4059 173 4059 173 4 b[24]
rlabel metal2 5139 177 5139 177 4 bb[22]
rlabel metal2 5351 177 5351 177 4 b[22]
rlabel metal2 6011 177 6011 177 4 bb[20]
rlabel metal2 6223 177 6223 177 4 b[20]
rlabel metal2 6883 177 6883 177 4 bb[18]
rlabel metal2 7095 177 7095 177 4 b[18]
rlabel metal2 7755 177 7755 177 4 bb[16]
rlabel metal2 7967 177 7967 177 4 b[16]
rlabel metal2 9045 175 9045 175 4 bb[14]
rlabel metal2 9257 175 9257 175 4 b[14]
rlabel metal2 9917 175 9917 175 4 bb[12]
rlabel metal2 10129 175 10129 175 4 b[12]
rlabel metal2 10789 175 10789 175 4 bb[10]
rlabel metal2 11001 175 11001 175 4 b[10]
rlabel metal2 11661 175 11661 175 4 bb[8]
rlabel metal2 11873 175 11873 175 4 b[8]
rlabel metal2 12957 181 12957 181 4 bb[6]
rlabel metal2 13169 181 13169 181 4 b[6]
rlabel metal2 13829 181 13829 181 4 bb[4]
rlabel metal2 14041 181 14041 181 4 b[4]
rlabel metal2 14701 181 14701 181 4 bb[2]
rlabel metal2 14913 181 14913 181 4 b[2]
rlabel metal2 15573 181 15573 181 4 bb[0]
rlabel metal2 15785 181 15785 181 4 b[0]
<< end >>
