magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nsubdiff >>
rect -36 49 36 62
rect -36 -49 -23 49
rect 23 -49 36 49
rect -36 -62 36 -49
<< nsubdiffcont >>
rect -23 -49 23 49
<< metal1 >>
rect -30 49 30 56
rect -30 -49 -23 49
rect 23 -49 30 49
rect -30 -56 30 -49
<< end >>
