magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< nwell >>
rect -174 -86 230 1356
<< pmos >>
rect 0 0 56 1270
<< pdiff >>
rect -88 1257 0 1270
rect -88 13 -75 1257
rect -29 13 0 1257
rect -88 0 0 13
rect 56 1257 144 1270
rect 56 13 85 1257
rect 131 13 144 1257
rect 56 0 144 13
<< pdiffc >>
rect -75 13 -29 1257
rect 85 13 131 1257
<< polysilicon >>
rect 0 1270 56 1314
rect 0 -44 56 0
<< metal1 >>
rect -75 1257 -29 1270
rect -75 0 -29 13
rect 85 1257 131 1270
rect 85 0 131 13
<< labels >>
flabel pdiffc -40 635 -40 635 0 FreeSans 186 0 0 0 S
flabel pdiffc 96 635 96 635 0 FreeSans 186 0 0 0 D
<< end >>
