magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal1 >>
rect -487 26 487 46
rect -487 -26 -469 26
rect 469 -26 487 26
rect -487 -46 487 -26
<< via1 >>
rect -469 -26 469 26
<< metal2 >>
rect -487 26 487 46
rect -487 -26 -469 26
rect 469 -26 487 26
rect -487 -46 487 -26
<< end >>
