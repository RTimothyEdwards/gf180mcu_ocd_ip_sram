magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal2 >>
rect -35 56 35 63
rect -35 -56 -28 56
rect 28 -56 35 56
rect -35 -63 35 -56
<< via2 >>
rect -28 -56 28 56
<< metal3 >>
rect -35 56 35 63
rect -35 -56 -28 56
rect 28 -56 35 56
rect -35 -63 35 -56
<< end >>
