magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal2 >>
rect -45 28 340 46
rect -45 -28 -28 28
rect 324 -28 340 28
rect -45 -46 340 -28
<< via2 >>
rect -28 -28 324 28
<< metal3 >>
rect -45 28 340 46
rect -45 -28 -28 28
rect 324 -28 340 28
rect -45 -46 340 -28
<< end >>
