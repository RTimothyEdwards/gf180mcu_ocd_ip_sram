magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< nwell >>
rect -194 -66 220 1483
<< polysilicon >>
rect -14 1418 41 1451
rect -14 -34 41 0
use pmos_5p04310591302067_3v512x8m81  pmos_5p04310591302067_3v512x8m81_0
timestamp 1763765945
transform 1 0 -14 0 1 0
box -174 -86 230 1504
<< end >>
