magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< error_s >>
rect 0 74 65 88
rect 0 17 3 74
rect 0 0 65 17
use via1_R90_512x8m81  via1_R90_512x8m81_0
timestamp 1763765945
transform 1 0 0 0 1 0
box 0 0 65 89
use via2_R90_512x8m81  via2_R90_512x8m81_0
timestamp 1763765945
transform 1 0 0 0 1 0
box 0 0 65 89
<< end >>
