magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -113 1148 113 1155
rect -113 -1148 -106 1148
rect 106 -1148 113 1148
rect -113 -1155 113 -1148
<< via2 >>
rect -106 -1148 106 1148
<< metal3 >>
rect -113 1148 113 1155
rect -113 -1148 -106 1148
rect 106 -1148 113 1148
rect -113 -1155 113 -1148
<< end >>
