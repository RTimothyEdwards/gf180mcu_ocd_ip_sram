magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal1 >>
rect -45 864 45 884
rect -45 -864 -26 864
rect 26 -864 45 864
rect -45 -884 45 -864
<< via1 >>
rect -26 -864 26 864
<< metal2 >>
rect -45 864 45 884
rect -45 -864 -26 864
rect 26 -864 45 864
rect -45 -884 45 -864
<< end >>
