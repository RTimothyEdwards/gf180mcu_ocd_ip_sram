magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal2 >>
rect -75 3376 45 7157
rect 150 3138 270 6934
rect 360 2900 480 6705
rect 570 2662 690 6482
rect 783 2424 903 6201
rect 994 2186 1114 5977
rect 1198 1948 1318 5740
rect 1425 1710 1545 5494
<< metal3 >>
rect -73 7038 1856 7189
rect 150 6793 1856 6944
rect 357 6548 1856 6699
rect 559 6303 1856 6453
rect 776 6082 1856 6232
rect 978 5839 1856 5990
rect 1174 5589 1856 5740
rect 1413 5345 1856 5496
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_0
timestamp 1763765945
transform -1 0 -7 0 1 3453
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_1
timestamp 1763765945
transform -1 0 219 0 1 3211
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_2
timestamp 1763765945
transform -1 0 429 0 1 2987
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_3
timestamp 1763765945
transform -1 0 640 0 1 2747
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_4
timestamp 1763765945
transform -1 0 853 0 1 2513
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_5
timestamp 1763765945
transform -1 0 1064 0 1 2252
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_6
timestamp 1763765945
transform -1 0 1268 0 1 2027
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_7
timestamp 1763765945
transform -1 0 1485 0 1 1790
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_8
timestamp 1763765945
transform -1 0 1268 0 1 5666
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_9
timestamp 1763765945
transform -1 0 1064 0 1 5916
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_10
timestamp 1763765945
transform -1 0 853 0 1 6158
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_11
timestamp 1763765945
transform -1 0 640 0 1 6379
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_12
timestamp 1763765945
transform -1 0 429 0 1 6624
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_13
timestamp 1763765945
transform -1 0 219 0 1 6865
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_14
timestamp 1763765945
transform -1 0 -7 0 1 7110
box -63 -63 63 63
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_15
timestamp 1763765945
transform -1 0 1492 0 1 5420
box -63 -63 63 63
<< end >>
