magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< polysilicon >>
rect -128 23 128 36
rect -128 -23 -114 23
rect 114 -23 128 23
rect -128 -36 128 -23
<< polycontact >>
rect -114 -23 114 23
<< metal1 >>
rect -122 23 122 30
rect -122 -23 -114 23
rect 114 -23 122 23
rect -122 -30 122 -23
<< end >>
