magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< nmos >>
rect 0 0 56 943
<< ndiff >>
rect -88 930 0 943
rect -88 13 -75 930
rect -29 13 0 930
rect -88 0 0 13
rect 56 930 144 943
rect 56 13 85 930
rect 131 13 144 930
rect 56 0 144 13
<< ndiffc >>
rect -75 13 -29 930
rect 85 13 131 930
<< polysilicon >>
rect 0 943 56 987
rect 0 -44 56 0
<< metal1 >>
rect -75 930 -29 943
rect -75 0 -29 13
rect 85 930 131 943
rect 85 0 131 13
<< labels >>
flabel ndiffc -40 471 -40 471 0 FreeSans 93 0 0 0 S
flabel ndiffc 96 471 96 471 0 FreeSans 93 0 0 0 D
<< end >>
