magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< error_p >>
rect -75 0 -29 84
rect 122 0 168 84
<< nwell >>
rect -174 -86 267 170
<< pmos >>
rect 0 0 93 84
<< pdiff >>
rect -88 71 0 84
rect -88 13 -75 71
rect -29 13 0 71
rect -88 0 0 13
rect 93 71 181 84
rect 93 13 122 71
rect 168 13 181 71
rect 93 0 181 13
<< pdiffc >>
rect -75 13 -29 71
rect 122 13 168 71
<< polysilicon >>
rect 0 84 93 128
rect 0 -44 93 0
<< metal1 >>
rect -75 71 -29 84
rect -75 0 -29 13
rect 122 71 168 84
rect 122 0 168 13
<< labels >>
flabel pdiffc -40 42 -40 42 0 FreeSans 186 0 0 0 S
flabel pdiffc 133 42 133 42 0 FreeSans 186 0 0 0 D
<< end >>
