magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal3 >>
rect 349 1275 1049 1701
use M2_M14310591302017_256x8m81  M2_M14310591302017_256x8m81_0
timestamp 1763564386
transform 1 0 699 0 1 1390
box -330 -113 330 113
use M3_M24310591302016_256x8m81  M3_M24310591302016_256x8m81_0
timestamp 1763564386
transform 1 0 699 0 1 1390
box -330 -113 330 113
<< end >>
