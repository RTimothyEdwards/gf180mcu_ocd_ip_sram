magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal1 >>
rect -8 189 75 215
rect -8 26 7 189
rect 59 26 75 189
rect -8 0 75 26
<< via1 >>
rect 7 26 59 189
<< metal2 >>
rect -8 189 75 215
rect -8 26 7 189
rect 59 26 75 189
rect -8 0 75 26
<< end >>
