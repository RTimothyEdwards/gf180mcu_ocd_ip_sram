magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< psubdiff >>
rect -970 71 970 109
rect -970 -71 -930 71
rect 930 -71 970 71
rect -970 -109 970 -71
<< psubdiffcont >>
rect -930 -71 930 71
<< metal1 >>
rect -956 71 956 95
rect -956 -71 -930 71
rect 930 -71 956 71
rect -956 -95 956 -71
<< end >>
