magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< nwell >>
rect -1758 -210 1759 210
<< nsubdiff >>
rect -1655 71 1655 109
rect -1655 -71 -1615 71
rect 1615 -71 1655 71
rect -1655 -109 1655 -71
<< nsubdiffcont >>
rect -1615 -71 1615 71
<< metal1 >>
rect -1641 71 1641 95
rect -1641 -71 -1615 71
rect 1615 -71 1641 71
rect -1641 -95 1641 -71
<< end >>
