magic
tech gf180mcuD
magscale 1 10
timestamp 1765212052
<< error_s >>
rect 467 4958 525 5019
<< nwell >>
rect 441 20127 4028 20391
rect 441 18837 3465 20127
rect 441 17060 4028 18837
rect 3849 17042 4028 17060
rect 225 13110 440 13973
rect 1585 6973 2050 7109
<< metal1 >>
rect 309 18913 373 18974
rect 308 12055 349 12122
rect 3740 8593 3806 8960
rect 1894 7447 1953 7663
rect 2391 6877 2534 6974
rect 1677 2149 1729 2223
rect 1842 2196 1918 2223
rect 1834 2067 1918 2196
rect 2342 2067 2426 2233
rect 316 -467 550 -415
<< metal2 >>
rect 281 18965 333 18991
rect 277 12088 334 18965
rect 431 12517 487 13882
rect 1288 12591 1344 13849
rect 2197 12591 2259 13866
rect 3101 12592 3164 13863
rect 3878 12444 3934 13852
rect 3544 12380 3934 12444
rect 1450 8700 1516 12125
rect 699 8595 1350 8652
rect 327 1792 392 7321
rect 581 6998 648 7659
rect 581 6934 809 6998
rect 742 5635 809 6934
rect 1294 6905 1350 8595
rect 1294 6848 1419 6905
rect 591 5566 809 5635
rect 591 2865 658 5566
rect 1055 5549 1121 5971
rect 1363 5754 1419 6848
rect 1579 6863 1645 12101
rect 1708 8700 1774 12125
rect 2963 7357 3028 7470
rect 3284 7436 3350 7470
rect 3284 7369 3535 7436
rect 2963 7289 3104 7357
rect 3469 7270 3535 7369
rect 1579 6806 1991 6863
rect 935 5462 1121 5549
rect 1310 5697 1419 5754
rect 935 4955 1001 5462
rect 915 4880 1001 4955
rect 591 2740 690 2865
rect 634 1797 690 2740
rect 915 2420 981 4880
rect 1310 2821 1366 5697
rect 1589 5007 1647 5616
rect 1924 5047 1991 6806
rect 3740 6237 3806 8678
rect 3740 6167 3826 6237
rect 3076 5651 3300 5745
rect 3760 5711 3826 6167
rect 3239 5432 3300 5651
rect 3587 5643 3826 5711
rect 3587 5432 3645 5643
rect 1495 4968 1647 5007
rect 1736 4991 1991 5047
rect 1736 4768 1802 4991
rect 1579 4683 1802 4768
rect 1579 3841 1645 4683
rect 915 2330 1011 2420
rect 945 1787 1011 2330
rect 1309 2204 1370 2821
rect 1309 2146 1430 2204
rect 1367 1777 1430 2146
rect 1367 1716 1452 1777
rect 1389 598 1452 1716
rect 1389 535 2159 598
rect 2096 213 2159 535
<< metal3 >>
rect 0 15758 351 17141
rect 263 12144 3861 12304
rect 3845 10038 4055 11944
rect 467 4958 525 5019
rect 222 4386 1617 4448
rect 3938 3704 4055 4657
rect 3945 1939 4055 2257
use din_3v512x8m81  din_3v512x8m81_0
timestamp 1764525316
transform 1 0 226 0 1 6408
box -156 560 1824 6415
use M1_NACTIVE4310591302024_3v512x8m81  M1_NACTIVE4310591302024_3v512x8m81_0
timestamp 1764525316
transform 1 0 3909 0 1 2090
box -38 -128 36 128
use M2_M1$$45012012_3v512x8m81  M2_M1$$45012012_3v512x8m81_0
timestamp 1764525316
transform 1 0 1767 0 1 12254
box -562 -46 562 46
use M2_M1$$45013036_3v512x8m81  M2_M1$$45013036_3v512x8m81_0
timestamp 1764525316
transform 1 0 2839 0 1 12254
box -266 -46 266 46
use M2_M1431059130200_3v512x8m81  M2_M1431059130200_3v512x8m81_0
timestamp 1764525316
transform 0 -1 3614 1 0 5373
box -63 -34 63 34
use M2_M1431059130200_3v512x8m81  M2_M1431059130200_3v512x8m81_1
timestamp 1764525316
transform 0 -1 3273 1 0 5373
box -63 -34 63 34
use M2_M1431059130208_3v512x8m81  M2_M1431059130208_3v512x8m81_0
timestamp 1764525316
transform 0 -1 642 1 0 1823
box -34 -63 34 63
use M2_M1431059130208_3v512x8m81  M2_M1431059130208_3v512x8m81_1
timestamp 1764525316
transform 1 0 2126 0 1 272
box -34 -63 34 63
use M2_M14310591302020_3v512x8m81  M2_M14310591302020_3v512x8m81_0
timestamp 1764525316
transform 1 0 299 0 1 18941
box -35 -56 35 55
use M2_M14310591302020_3v512x8m81  M2_M14310591302020_3v512x8m81_1
timestamp 1764525316
transform 1 0 461 0 1 13884
box -35 -56 35 55
use M2_M14310591302020_3v512x8m81  M2_M14310591302020_3v512x8m81_2
timestamp 1764525316
transform 1 0 3901 0 1 13869
box -35 -56 35 55
use M2_M14310591302020_3v512x8m81  M2_M14310591302020_3v512x8m81_3
timestamp 1764525316
transform 1 0 307 0 1 12088
box -35 -56 35 55
use M2_M14310591302025_3v512x8m81  M2_M14310591302025_3v512x8m81_0
timestamp 1764525316
transform 1 0 3909 0 1 2091
box -34 -85 34 135
use m2_saout01_3v512x8m81  m2_saout01_3v512x8m81_0
timestamp 1764525316
transform 1 0 480 0 1 20290
box -102 -44 3491 1507
use M3_M2$$43370540_3v512x8m81  M3_M2$$43370540_3v512x8m81_0
timestamp 1764525316
transform 1 0 2839 0 1 12254
box -266 -46 266 46
use M3_M2$$44741676_3v512x8m81  M3_M2$$44741676_3v512x8m81_0
timestamp 1764525316
transform 1 0 1767 0 1 12254
box -562 -46 562 46
use M3_M2431059130207_3v512x8m81  M3_M2431059130207_3v512x8m81_0
timestamp 1764525316
transform 1 0 1554 0 1 4987
box -63 -35 63 35
use M3_M24310591302026_3v512x8m81  M3_M24310591302026_3v512x8m81_0
timestamp 1764525316
transform 1 0 3909 0 1 2091
box -35 -135 35 135
use mux821_3v512x8m81  mux821_3v512x8m81_0
timestamp 1765212052
transform 1 0 387 0 1 12008
box -575 634 4956 8484
use outbuf_oe_3v512x8m81  outbuf_oe_3v512x8m81_0
timestamp 1764693003
transform 1 0 442 0 1 5371
box -372 -251 3623 2214
use sa_3v512x8m81  sa_3v512x8m81_0
timestamp 1764525316
transform 1 0 442 0 1 6970
box -249 376 3523 5747
use sacntl_2_3v512x8m81  sacntl_2_3v512x8m81_0
timestamp 1764692725
transform 1 0 442 0 1 1531
box -371 244 3623 3958
use via1_2_x2_3v512x8m81  via1_2_x2_3v512x8m81_0
timestamp 1764525316
transform 1 0 1451 0 1 9585
box -9 0 73 215
use via1_2_x2_3v512x8m81  via1_2_x2_3v512x8m81_1
timestamp 1764525316
transform 1 0 1451 0 1 9222
box -9 0 73 215
use via1_2_x2_3v512x8m81  via1_2_x2_3v512x8m81_2
timestamp 1764525316
transform 1 0 1451 0 1 8901
box -9 0 73 215
use via1_x2_3v512x8m81  via1_x2_3v512x8m81_0
timestamp 1764525316
transform -1 0 1644 0 -1 12123
box -8 0 72 222
use via1_x2_3v512x8m81  via1_x2_3v512x8m81_1
timestamp 1764525316
transform -1 0 1122 0 -1 5966
box -8 0 72 222
use via1_x2_3v512x8m81  via1_x2_3v512x8m81_2
timestamp 1764525316
transform 1 0 1579 0 1 3842
box -8 0 72 222
use via1_x2_3v512x8m81  via1_x2_3v512x8m81_3
timestamp 1764525316
transform 1 0 3741 0 1 8517
box -8 0 72 222
use via1_x2_3v512x8m81  via1_x2_3v512x8m81_4
timestamp 1764525316
transform 1 0 322 0 1 7236
box -8 0 72 222
use via1_x2_R90_3v512x8m81  via1_x2_R90_3v512x8m81_0
timestamp 1764525316
transform 0 -1 3592 1 0 12378
box -8 0 72 215
use via1_x2_R90_3v512x8m81  via1_x2_R90_3v512x8m81_1
timestamp 1764525316
transform 0 -1 1381 1 0 13836
box -8 0 72 215
use via1_x2_R90_3v512x8m81  via1_x2_R90_3v512x8m81_2
timestamp 1764525316
transform 0 -1 2271 1 0 13836
box -8 0 72 215
use via1_x2_R90_3v512x8m81  via1_x2_R90_3v512x8m81_3
timestamp 1764525316
transform 0 -1 3185 1 0 13836
box -8 0 72 215
use via1_x2_R90_3v512x8m81  via1_x2_R90_3v512x8m81_4
timestamp 1764525316
transform 0 -1 647 1 0 7628
box -8 0 72 215
use via2_3v512x8m81  via2_3v512x8m81_0
timestamp 1764525316
transform 1 0 3743 0 1 13851
box 0 0 65 92
use via2_3v512x8m81  via2_3v512x8m81_1
timestamp 1764525316
transform 1 0 3135 0 1 14092
box 0 0 65 92
use via2_3v512x8m81  via2_3v512x8m81_2
timestamp 1764525316
transform 1 0 2947 0 1 14330
box 0 0 65 92
use via2_3v512x8m81  via2_3v512x8m81_3
timestamp 1764525316
transform 1 0 2046 0 1 14805
box 0 0 65 92
use via2_3v512x8m81  via2_3v512x8m81_4
timestamp 1764525316
transform 1 0 2229 0 1 14579
box 0 0 65 92
use via2_3v512x8m81  via2_3v512x8m81_5
timestamp 1764525316
transform 1 0 1331 0 1 15050
box 0 0 65 92
use via2_3v512x8m81  via2_3v512x8m81_6
timestamp 1764525316
transform 1 0 1143 0 1 15291
box 0 0 65 92
use via2_3v512x8m81  via2_3v512x8m81_7
timestamp 1764525316
transform 0 1 398 -1 0 15578
box 0 0 65 92
use via2_x2_3v512x8m81  via2_x2_3v512x8m81_0
timestamp 1764525316
transform 1 0 1709 0 1 9222
box -9 0 74 222
use via2_x2_3v512x8m81  via2_x2_3v512x8m81_1
timestamp 1764525316
transform 1 0 1709 0 1 9222
box -9 0 74 222
use via2_x2_3v512x8m81  via2_x2_3v512x8m81_2
timestamp 1764525316
transform 1 0 1709 0 1 9222
box -9 0 74 222
use via2_x2_3v512x8m81  via2_x2_3v512x8m81_3
timestamp 1764525316
transform 1 0 1709 0 1 9222
box -9 0 74 222
use via2_x2_3v512x8m81  via2_x2_3v512x8m81_4
timestamp 1764525316
transform 1 0 1709 0 1 8901
box -9 0 74 222
use via2_x2_3v512x8m81  via2_x2_3v512x8m81_5
timestamp 1764525316
transform 1 0 1709 0 1 9585
box -9 0 74 222
use wen_wm1_3v512x8m81  wen_wm1_3v512x8m81_0
timestamp 1764692000
transform 1 0 225 0 1 -451
box -139 -24 3471 2300
<< labels >>
rlabel metal3 s 653 20231 653 20231 4 vdd
port 10 nsew
rlabel metal2 s 3403 20112 3403 20112 4 bb[1]
port 16 nsew
rlabel metal2 s 2682 20115 2682 20115 4 bb[2]
port 18 nsew
rlabel metal2 s 2542 20118 2542 20118 4 bb[3]
port 19 nsew
rlabel metal2 s 1815 20113 1815 20113 4 bb[4]
port 20 nsew
rlabel metal2 s 1670 20113 1670 20113 4 bb[5]
port 21 nsew
rlabel metal2 s 808 20118 808 20118 4 bb[7]
port 22 nsew
rlabel metal2 s 948 20113 948 20113 4 bb[6]
port 23 nsew
rlabel metal2 s 3114 20112 3114 20112 4 b[1]
port 25 nsew
rlabel metal2 s 2104 20112 2104 20112 4 b[4]
port 26 nsew
rlabel metal2 s 1380 20112 1380 20112 4 b[5]
port 27 nsew
rlabel metal2 s 1239 20112 1239 20112 4 b[6]
port 28 nsew
rlabel metal2 s 515 20112 515 20112 4 b[7]
port 29 nsew
rlabel metal2 s 2975 20112 2975 20112 4 b[2]
port 30 nsew
rlabel metal2 s 2247 20112 2247 20112 4 b[3]
port 31 nsew
rlabel metal2 s 511 20112 511 20112 4 b[7]
port 29 nsew
rlabel metal2 s 1237 20112 1237 20112 4 b[6]
port 28 nsew
rlabel metal2 s 1383 20112 1383 20112 4 b[5]
port 27 nsew
rlabel metal2 s 2102 20112 2102 20112 4 b[4]
port 26 nsew
rlabel metal2 s 2245 20112 2245 20112 4 b[3]
port 31 nsew
rlabel metal2 s 2974 20112 2974 20112 4 b[2]
port 30 nsew
rlabel metal2 s 3115 20112 3115 20112 4 b[1]
port 25 nsew
rlabel metal2 s 947 20113 947 20113 4 bb[6]
port 23 nsew
rlabel metal2 s 805 20118 805 20118 4 bb[7]
port 22 nsew
rlabel metal2 s 1673 20113 1673 20113 4 bb[5]
port 21 nsew
rlabel metal2 s 1813 20113 1813 20113 4 bb[4]
port 20 nsew
rlabel metal2 s 2539 20118 2539 20118 4 bb[3]
port 19 nsew
rlabel metal2 s 2679 20115 2679 20115 4 bb[2]
port 18 nsew
rlabel metal2 s 3404 20112 3404 20112 4 bb[1]
port 16 nsew
rlabel metal3 s 567 14482 567 14482 4 ypass[4]
port 4 nsew
rlabel metal3 s 567 15153 567 15153 4 ypass[7]
port 7 nsew
rlabel metal3 s 567 14931 567 14931 4 ypass[6]
port 6 nsew
rlabel metal3 s 567 14709 567 14709 4 ypass[5]
port 5 nsew
rlabel metal3 s 567 14023 567 14023 4 ypass[3]
port 3 nsew
rlabel metal3 s 567 13801 567 13801 4 ypass[2]
port 2 nsew
rlabel metal3 s 567 13579 567 13579 4 ypass[1]
port 1 nsew
rlabel metal3 s 664 15750 664 15750 4 vss
port 9 nsew
rlabel metal3 s 567 13354 567 13354 4 ypass[0]
port 11 nsew
rlabel metal1 s 695 19297 695 19297 4 pcb
port 34 nsew
rlabel metal1 s 695 19295 695 19295 4 pcb
port 34 nsew
flabel metal3 s 322 16817 322 16817 0 FreeSans 420 0 0 0 VSS
port 14 nsew
rlabel metal1 s 1260 12099 1260 12099 4 pcb
port 34 nsew
rlabel metal1 s 488 6764 488 6764 4 datain
port 32 nsew
flabel metal3 s 322 10195 322 10195 0 FreeSans 420 0 0 0 VDD
port 12 nsew
flabel metal3 s 322 6915 322 6915 0 FreeSans 420 0 0 0 VDD
port 12 nsew
flabel metal3 s 322 9710 322 9710 0 FreeSans 420 0 0 0 VSS
port 14 nsew
rlabel metal3 s 1264 10577 1264 10577 4 vdd
port 10 nsew
rlabel metal3 s 681 12768 681 12768 4 vss
port 9 nsew
rlabel metal3 s 1314 8665 1314 8665 4 vss
port 9 nsew
flabel metal3 s 449 13455 449 13455 0 FreeSans 420 0 0 0 VDD
port 12 nsew
flabel metal3 s 453 12893 453 12893 0 FreeSans 420 0 0 0 VSS
port 14 nsew
rlabel metal3 s 616 2536 616 2536 4 men
port 8 nsew
rlabel metal3 s 2121 4191 2121 4191 4 vdd
port 10 nsew
rlabel metal3 s 1484 1794 1484 1794 4 vdd
port 10 nsew
rlabel metal3 s 1957 5339 1957 5339 4 vss
port 9 nsew
rlabel metal3 s 2312 6862 2312 6862 4 vdd
port 10 nsew
flabel metal3 s 322 6478 322 6478 0 FreeSans 420 0 0 0 VDD
port 12 nsew
flabel metal3 s 322 3826 322 3826 0 FreeSans 420 0 0 0 VDD
port 12 nsew
flabel metal3 s 322 3238 322 3238 0 FreeSans 420 0 0 0 VSS
port 14 nsew
flabel metal3 s 322 5938 322 5938 0 FreeSans 420 0 0 0 VSS
port 14 nsew
rlabel metal2 s 975 2301 975 2301 4 q
port 33 nsew
rlabel metal2 s 346 2721 346 2721 4 datain
port 32 nsew
flabel metal3 s 322 1497 322 1497 0 FreeSans 420 0 0 0 VDD
port 12 nsew
flabel metal3 s 322 -133 322 -133 0 FreeSans 420 0 0 0 VDD
port 12 nsew
flabel metal3 s 431 508 431 508 0 FreeSans 420 0 0 0 GWEN
port 13 nsew
flabel metal3 s 322 336 322 336 0 FreeSans 420 0 0 0 VSS
port 14 nsew
flabel metal3 s 322 981 322 981 0 FreeSans 420 0 0 0 VSS
port 14 nsew
flabel metal3 s 322 671 322 671 0 FreeSans 420 0 0 0 VSS
port 14 nsew
flabel metal1 s 505 -443 505 -443 0 FreeSans 420 0 0 0 WEN
port 35 nsew
flabel metal3 s 322 2466 322 2466 0 FreeSans 420 0 0 0 VSS
port 14 nsew
flabel metal3 s 322 2125 322 2125 0 FreeSans 420 0 0 0 VDD
port 12 nsew
rlabel metal3 s 2042 2573 2042 2573 4 vss
port 9 nsew
rlabel metal3 s 2042 3235 2042 3235 4 vss
port 9 nsew
rlabel metal3 s 653 13454 653 13454 4 vdd
port 10 nsew
flabel metal3 s 480 4986 480 4986 0 FreeSans 420 0 0 0 GWE
port 15 nsew
<< end >>
