magic
tech gf180mcuD
magscale 1 10
timestamp 1765833244
<< metal2 >>
rect -782 28 783 46
rect -782 -28 -766 28
rect 766 -28 783 28
rect -782 -46 783 -28
<< via2 >>
rect -766 -28 766 28
<< metal3 >>
rect -783 28 783 46
rect -783 -28 -766 28
rect 766 -28 783 28
rect -783 -46 783 -28
<< end >>
