magic
tech gf180mcuD
magscale 1 10
timestamp 1765833244
<< psubdiff >>
rect -56 169 56 203
rect -56 -709 -23 169
rect 23 -709 56 169
rect -56 -742 56 -709
<< psubdiffcont >>
rect -23 -709 23 169
<< metal1 >>
rect -49 169 49 197
rect -49 -709 -23 169
rect 23 -709 49 169
rect -49 -737 49 -709
<< end >>
