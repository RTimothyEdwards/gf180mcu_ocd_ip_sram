magic
tech gf180mcuD
magscale 1 10
timestamp 1763564386
<< metal2 >>
rect -118 333 119 351
rect -118 -333 -102 333
rect 102 -333 119 333
rect -118 -351 119 -333
<< via2 >>
rect -102 -333 102 333
<< metal3 >>
rect -119 333 119 351
rect -119 -333 -102 333
rect 102 -333 119 333
rect -119 -351 119 -333
<< end >>
