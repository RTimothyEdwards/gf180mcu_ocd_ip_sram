magic
tech gf180mcuD
magscale 1 10
timestamp 1763477050
<< metal2 >>
rect -4 1821 151 13188
rect 346 2486 503 11480
rect 707 1821 863 13180
use M2_M14310591302097_512x8m81  M2_M14310591302097_512x8m81_0
timestamp 1763476864
transform 1 0 784 0 1 2160
box -70 -330 70 330
use M2_M14310591302097_512x8m81  M2_M14310591302097_512x8m81_1
timestamp 1763476864
transform 1 0 72 0 1 2160
box -70 -330 70 330
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_0
timestamp 1763476864
transform 1 0 424 0 1 4635
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_1
timestamp 1763476864
transform 1 0 786 0 1 3508
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_2
timestamp 1763476864
transform 1 0 74 0 1 4157
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_3
timestamp 1763476864
transform 1 0 786 0 1 4157
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_4
timestamp 1763476864
transform 1 0 424 0 1 5389
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_5
timestamp 1763476864
transform 1 0 786 0 1 5808
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_6
timestamp 1763476864
transform 1 0 74 0 1 5808
box -70 -113 70 113
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_7
timestamp 1763476864
transform 1 0 74 0 1 3508
box -70 -113 70 113
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_0
timestamp 1763476864
transform 1 0 74 0 1 6728
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_1
timestamp 1763476864
transform 1 0 74 0 1 9451
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_2
timestamp 1763476864
transform 1 0 786 0 1 9451
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_3
timestamp 1763476864
transform 1 0 74 0 1 8970
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_4
timestamp 1763476864
transform 1 0 786 0 1 8970
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_5
timestamp 1763476864
transform 1 0 74 0 1 12935
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_6
timestamp 1763476864
transform 1 0 786 0 1 12935
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_7
timestamp 1763476864
transform 1 0 74 0 1 12454
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_8
timestamp 1763476864
transform 1 0 786 0 1 12454
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_9
timestamp 1763476864
transform 1 0 74 0 1 11975
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_10
timestamp 1763476864
transform 1 0 786 0 1 11975
box -70 -200 70 200
use M3_M24310591302098_512x8m81  M3_M24310591302098_512x8m81_11
timestamp 1763476864
transform 1 0 786 0 1 6728
box -70 -200 70 200
use M3_M24310591302099_512x8m81  M3_M24310591302099_512x8m81_0
timestamp 1763476864
transform 1 0 424 0 1 10800
box -70 -634 70 634
use M3_M243105913020100_512x8m81  M3_M243105913020100_512x8m81_0
timestamp 1763476864
transform 1 0 424 0 1 7792
box -70 -417 70 417
use M3_M243105913020101_512x8m81  M3_M243105913020101_512x8m81_0
timestamp 1763476864
transform 1 0 424 0 1 2843
box -70 -330 70 330
<< end >>
