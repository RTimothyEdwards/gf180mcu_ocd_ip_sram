magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_0
timestamp 1763766357
transform -1 0 7817 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_1
timestamp 1763766357
transform -1 0 8689 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_2
timestamp 1763766357
transform -1 0 8253 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_3
timestamp 1763766357
transform -1 0 9125 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_4
timestamp 1763766357
transform -1 0 9561 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_5
timestamp 1763766357
transform -1 0 9997 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_6
timestamp 1763766357
transform -1 0 10433 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_7
timestamp 1763766357
transform -1 0 6525 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_8
timestamp 1763766357
transform -1 0 6089 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_9
timestamp 1763766357
transform -1 0 5653 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_10
timestamp 1763766357
transform -1 0 5217 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_11
timestamp 1763766357
transform -1 0 4345 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_12
timestamp 1763766357
transform -1 0 4781 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_13
timestamp 1763766357
transform -1 0 3909 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_14
timestamp 1763766357
transform -1 0 3473 0 1 177
box 62 89 538 797
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_15
timestamp 1763766357
transform -1 0 7381 0 1 177
box 62 89 538 797
use 018SRAM_strap1_256x8m81  018SRAM_strap1_256x8m81_0
timestamp 1763766357
transform -1 0 6954 0 1 177
box 91 55 511 797
use 018SRAM_strap1_256x8m81  018SRAM_strap1_256x8m81_1
timestamp 1763766357
transform -1 0 10862 0 1 177
box 91 55 511 797
<< end >>
