magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< polysilicon >>
rect -14 635 41 669
rect -14 -34 41 0
use nmos_5p0431059130200_3v1024x8m81  nmos_5p0431059130200_3v1024x8m81_0
timestamp 1764525316
transform 1 0 -14 0 1 0
box -88 -44 144 679
<< end >>
