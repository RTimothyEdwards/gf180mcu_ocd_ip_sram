magic
tech gf180mcuD
magscale 1 10
timestamp 1764700137
<< psubdiff >>
rect -165 73 166 114
rect -165 -73 -126 73
rect 126 -73 166 73
rect -165 -114 166 -73
<< psubdiffcont >>
rect -126 -73 126 73
<< metal1 >>
rect -159 73 160 108
rect -159 -73 -126 73
rect 126 -73 160 73
rect -159 -107 160 -73
<< end >>
