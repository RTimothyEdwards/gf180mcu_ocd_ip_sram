magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect -174 -86 230 721
<< pmos >>
rect 0 0 56 635
<< pdiff >>
rect -88 622 0 635
rect -88 13 -75 622
rect -29 13 0 622
rect -88 0 0 13
rect 56 622 144 635
rect 56 13 85 622
rect 131 13 144 622
rect 56 0 144 13
<< pdiffc >>
rect -75 13 -29 622
rect 85 13 131 622
<< polysilicon >>
rect 0 635 56 679
rect 0 -44 56 0
<< metal1 >>
rect -75 622 -29 635
rect -75 0 -29 13
rect 85 622 131 635
rect 85 0 131 13
<< labels >>
flabel pdiffc -40 317 -40 317 0 FreeSans 186 0 0 0 S
flabel pdiffc 96 317 96 317 0 FreeSans 186 0 0 0 D
<< end >>
