magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect -154 -1302 154 1302
<< nsubdiff >>
rect -54 1166 53 1199
rect -54 -1166 -23 1166
rect 23 -1166 53 1166
rect -54 -1198 53 -1166
<< nsubdiffcont >>
rect -23 -1166 23 1166
<< metal1 >>
rect -40 1166 40 1184
rect -40 -1166 -23 1166
rect 23 -1166 40 1166
rect -40 -1184 40 -1166
<< end >>
