VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_ocd_ip_sram__sram512x8m8wm1
  CLASS BLOCK ;
  FOREIGN gf180mcu_ocd_ip_sram__sram512x8m8wm1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 301.300 BY 321.890 ;
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 101.520 0.000 102.305 6.000 ;
    END
  END A[8]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 103.965 0.000 104.750 6.000 ;
    END
  END A[7]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 188.200 0.000 188.985 6.000 ;
    END
  END A[6]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 190.455 0.000 191.240 6.000 ;
    END
  END A[5]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 193.070 0.000 193.855 6.000 ;
    END
  END A[4]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 196.925 0.000 197.710 6.000 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 108.005 0.000 108.790 6.000 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 113.930 0.000 114.715 6.000 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 119.850 0.000 120.630 6.000 ;
    END
  END A[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.928400 ;
    PORT
      LAYER Metal2 ;
        RECT 176.195 0.000 176.980 6.000 ;
    END
  END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.738400 ;
    PORT
      LAYER Metal2 ;
        RECT 97.775 0.000 98.560 6.000 ;
    END
  END CLK
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 291.200 5.030 291.985 6.000 ;
        RECT 290.800 4.305 291.985 5.030 ;
        RECT 290.800 0.000 291.585 4.305 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 254.645 4.245 254.930 6.000 ;
        RECT 254.605 0.000 255.385 4.245 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 249.530 4.245 249.810 6.000 ;
        RECT 249.235 0.000 250.020 4.245 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 212.255 4.355 212.625 6.000 ;
        RECT 212.255 4.350 213.940 4.355 ;
        RECT 212.255 3.985 214.845 4.350 ;
        RECT 214.060 0.000 214.845 3.985 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 85.695 4.850 86.000 6.000 ;
        RECT 83.280 4.545 86.000 4.850 ;
        RECT 83.280 0.000 84.065 4.545 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 48.730 5.425 49.015 6.000 ;
        RECT 47.595 5.140 49.015 5.425 ;
        RECT 47.595 4.160 47.880 5.140 ;
        RECT 47.085 3.720 47.880 4.160 ;
        RECT 47.085 0.000 47.870 3.720 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 43.215 5.290 43.540 6.000 ;
        RECT 43.180 4.170 43.540 5.290 ;
        RECT 42.720 0.000 43.505 4.170 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.249200 ;
    PORT
      LAYER Metal2 ;
        RECT 6.520 0.000 7.305 6.000 ;
    END
  END D[0]
  PIN GWEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.141600 ;
    PORT
      LAYER Metal2 ;
        RECT 142.055 0.000 142.840 6.000 ;
    END
  END GWEN
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 285.870 4.245 286.200 6.000 ;
        RECT 285.490 0.000 286.275 4.245 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 257.025 4.245 257.345 6.000 ;
        RECT 256.960 0.000 257.740 4.245 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 247.175 4.245 247.460 6.000 ;
        RECT 246.880 0.000 247.665 4.245 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 217.860 4.705 218.190 6.000 ;
        RECT 217.860 4.695 220.060 4.705 ;
        RECT 217.860 4.375 220.135 4.695 ;
        RECT 219.350 0.000 220.135 4.375 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 77.980 4.130 78.315 6.000 ;
        RECT 77.975 0.000 78.760 4.130 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 51.250 5.450 51.580 6.000 ;
        RECT 49.960 5.120 51.580 5.450 ;
        RECT 49.960 4.160 50.290 5.120 ;
        RECT 49.440 3.710 50.290 4.160 ;
        RECT 49.440 0.000 50.225 3.710 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 41.545 4.725 41.875 6.000 ;
        RECT 40.840 4.395 41.875 4.725 ;
        RECT 40.840 4.200 41.170 4.395 ;
        RECT 40.365 3.555 41.170 4.200 ;
        RECT 40.365 0.000 41.145 3.555 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.315450 ;
    PORT
      LAYER Metal2 ;
        RECT 12.255 5.780 12.585 6.000 ;
        RECT 12.255 5.450 14.415 5.780 ;
        RECT 14.085 4.245 14.415 5.450 ;
        RECT 13.830 0.000 14.610 4.245 ;
    END
  END Q[0]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT 103.900 315.890 194.020 316.770 ;
        RECT 7.680 5.780 25.360 6.000 ;
        RECT 29.080 5.780 64.190 6.000 ;
        RECT 29.080 5.770 46.760 5.780 ;
        RECT 67.910 5.770 85.590 6.000 ;
        RECT 212.985 5.780 230.665 6.000 ;
        RECT 234.385 5.785 269.745 6.000 ;
        RECT 234.385 5.770 252.065 5.785 ;
        RECT 273.465 5.775 291.145 6.000 ;
      LAYER Metal1 ;
        RECT 4.845 311.335 5.975 312.050 ;
        RECT 4.845 310.635 6.000 311.335 ;
        RECT 295.440 311.080 296.570 312.135 ;
        RECT 295.300 310.800 296.570 311.080 ;
        RECT 4.845 309.620 5.975 310.635 ;
        RECT 295.440 309.705 296.570 310.800 ;
        RECT 4.845 305.275 5.975 305.990 ;
        RECT 4.845 304.575 6.000 305.275 ;
        RECT 295.440 305.020 296.570 306.075 ;
        RECT 295.300 304.740 296.570 305.020 ;
        RECT 4.845 303.560 5.975 304.575 ;
        RECT 295.440 303.645 296.570 304.740 ;
        RECT 4.845 299.215 5.975 299.930 ;
        RECT 4.845 298.515 6.000 299.215 ;
        RECT 295.440 298.960 296.570 300.015 ;
        RECT 295.300 298.680 296.570 298.960 ;
        RECT 4.845 297.500 5.975 298.515 ;
        RECT 295.440 297.585 296.570 298.680 ;
        RECT 4.845 293.155 5.975 293.870 ;
        RECT 4.845 292.455 6.000 293.155 ;
        RECT 295.440 292.900 296.570 293.955 ;
        RECT 295.300 292.620 296.570 292.900 ;
        RECT 4.845 291.440 5.975 292.455 ;
        RECT 295.440 291.525 296.570 292.620 ;
        RECT 4.845 287.095 5.975 287.810 ;
        RECT 4.845 286.395 6.000 287.095 ;
        RECT 295.440 286.840 296.570 287.895 ;
        RECT 295.300 286.560 296.570 286.840 ;
        RECT 4.845 285.380 5.975 286.395 ;
        RECT 295.440 285.465 296.570 286.560 ;
        RECT 4.845 281.035 5.975 281.750 ;
        RECT 4.845 280.335 6.000 281.035 ;
        RECT 295.440 280.780 296.570 281.835 ;
        RECT 295.300 280.500 296.570 280.780 ;
        RECT 4.845 279.320 5.975 280.335 ;
        RECT 295.440 279.405 296.570 280.500 ;
        RECT 4.845 274.975 5.975 275.690 ;
        RECT 4.845 274.275 6.000 274.975 ;
        RECT 295.440 274.720 296.570 275.775 ;
        RECT 295.300 274.440 296.570 274.720 ;
        RECT 4.845 273.260 5.975 274.275 ;
        RECT 295.440 273.345 296.570 274.440 ;
        RECT 4.845 268.915 5.975 269.630 ;
        RECT 4.845 268.215 6.000 268.915 ;
        RECT 295.440 268.660 296.570 269.715 ;
        RECT 295.300 268.380 296.570 268.660 ;
        RECT 4.845 267.200 5.975 268.215 ;
        RECT 295.440 267.285 296.570 268.380 ;
        RECT 4.845 262.855 5.975 263.570 ;
        RECT 4.845 262.155 6.000 262.855 ;
        RECT 295.440 262.600 296.570 263.655 ;
        RECT 295.300 262.320 296.570 262.600 ;
        RECT 4.845 261.140 5.975 262.155 ;
        RECT 295.440 261.225 296.570 262.320 ;
        RECT 4.845 256.795 5.975 257.510 ;
        RECT 4.845 256.095 6.000 256.795 ;
        RECT 295.440 256.540 296.570 257.595 ;
        RECT 295.300 256.260 296.570 256.540 ;
        RECT 4.845 255.080 5.975 256.095 ;
        RECT 295.440 255.165 296.570 256.260 ;
        RECT 4.845 250.735 5.975 251.450 ;
        RECT 4.845 250.035 6.000 250.735 ;
        RECT 295.440 250.480 296.570 251.535 ;
        RECT 295.300 250.200 296.570 250.480 ;
        RECT 4.845 249.020 5.975 250.035 ;
        RECT 295.440 249.105 296.570 250.200 ;
        RECT 4.845 244.675 5.975 245.390 ;
        RECT 4.845 243.975 6.000 244.675 ;
        RECT 295.440 244.420 296.570 245.475 ;
        RECT 295.300 244.140 296.570 244.420 ;
        RECT 4.845 242.960 5.975 243.975 ;
        RECT 295.440 243.045 296.570 244.140 ;
        RECT 4.845 238.615 5.975 239.330 ;
        RECT 4.845 237.915 6.000 238.615 ;
        RECT 295.440 238.360 296.570 239.415 ;
        RECT 295.300 238.080 296.570 238.360 ;
        RECT 4.845 236.900 5.975 237.915 ;
        RECT 295.440 236.985 296.570 238.080 ;
        RECT 4.845 232.555 5.975 233.270 ;
        RECT 4.845 231.855 6.000 232.555 ;
        RECT 295.440 232.300 296.570 233.355 ;
        RECT 295.300 232.020 296.570 232.300 ;
        RECT 4.845 230.840 5.975 231.855 ;
        RECT 295.440 230.925 296.570 232.020 ;
        RECT 4.845 226.495 5.975 227.210 ;
        RECT 4.845 225.795 6.000 226.495 ;
        RECT 295.440 226.240 296.570 227.295 ;
        RECT 295.300 225.960 296.570 226.240 ;
        RECT 4.845 224.780 5.975 225.795 ;
        RECT 295.440 224.865 296.570 225.960 ;
        RECT 4.845 220.435 5.975 221.150 ;
        RECT 4.845 219.735 6.000 220.435 ;
        RECT 295.440 220.180 296.570 221.235 ;
        RECT 295.300 219.900 296.570 220.180 ;
        RECT 4.845 218.720 5.975 219.735 ;
        RECT 295.440 218.805 296.570 219.900 ;
        RECT 4.845 214.375 5.975 215.090 ;
        RECT 4.845 213.675 6.000 214.375 ;
        RECT 295.440 214.120 296.570 215.175 ;
        RECT 295.300 213.840 296.570 214.120 ;
        RECT 4.845 212.660 5.975 213.675 ;
        RECT 295.440 212.745 296.570 213.840 ;
        RECT 4.845 208.315 5.975 209.030 ;
        RECT 4.845 207.615 6.000 208.315 ;
        RECT 295.440 208.060 296.570 209.115 ;
        RECT 295.300 207.780 296.570 208.060 ;
        RECT 4.845 206.600 5.975 207.615 ;
        RECT 295.440 206.685 296.570 207.780 ;
        RECT 4.845 202.255 5.975 202.970 ;
        RECT 4.845 201.555 6.000 202.255 ;
        RECT 295.440 202.000 296.570 203.055 ;
        RECT 295.300 201.720 296.570 202.000 ;
        RECT 4.845 200.540 5.975 201.555 ;
        RECT 295.440 200.625 296.570 201.720 ;
        RECT 4.845 196.195 5.975 196.910 ;
        RECT 4.845 195.495 6.000 196.195 ;
        RECT 295.440 195.940 296.570 196.995 ;
        RECT 295.300 195.660 296.570 195.940 ;
        RECT 4.845 194.480 5.975 195.495 ;
        RECT 295.440 194.565 296.570 195.660 ;
        RECT 4.845 190.135 5.975 190.850 ;
        RECT 4.845 189.435 6.000 190.135 ;
        RECT 295.440 189.880 296.570 190.935 ;
        RECT 295.300 189.600 296.570 189.880 ;
        RECT 4.845 188.420 5.975 189.435 ;
        RECT 295.440 188.505 296.570 189.600 ;
        RECT 4.845 184.075 5.975 184.790 ;
        RECT 4.845 183.375 6.000 184.075 ;
        RECT 295.440 183.820 296.570 184.875 ;
        RECT 295.300 183.540 296.570 183.820 ;
        RECT 4.845 182.360 5.975 183.375 ;
        RECT 295.440 182.445 296.570 183.540 ;
        RECT 4.845 178.015 5.975 178.730 ;
        RECT 4.845 177.315 6.000 178.015 ;
        RECT 295.440 177.760 296.570 178.815 ;
        RECT 295.300 177.480 296.570 177.760 ;
        RECT 4.845 176.300 5.975 177.315 ;
        RECT 295.440 176.385 296.570 177.480 ;
        RECT 4.845 171.955 5.975 172.670 ;
        RECT 4.845 171.255 6.000 171.955 ;
        RECT 295.440 171.700 296.570 172.755 ;
        RECT 295.300 171.420 296.570 171.700 ;
        RECT 4.845 170.240 5.975 171.255 ;
        RECT 295.440 170.325 296.570 171.420 ;
        RECT 4.845 165.895 5.975 166.610 ;
        RECT 4.845 165.195 6.000 165.895 ;
        RECT 295.440 165.640 296.570 166.695 ;
        RECT 295.300 165.360 296.570 165.640 ;
        RECT 4.845 164.180 5.975 165.195 ;
        RECT 295.440 164.265 296.570 165.360 ;
        RECT 4.845 159.835 5.975 160.550 ;
        RECT 4.845 159.135 6.000 159.835 ;
        RECT 295.440 159.580 296.570 160.635 ;
        RECT 295.300 159.300 296.570 159.580 ;
        RECT 4.845 158.120 5.975 159.135 ;
        RECT 295.440 158.205 296.570 159.300 ;
        RECT 4.845 153.775 5.975 154.490 ;
        RECT 4.845 153.075 6.000 153.775 ;
        RECT 295.440 153.520 296.570 154.575 ;
        RECT 295.300 153.240 296.570 153.520 ;
        RECT 4.845 152.060 5.975 153.075 ;
        RECT 295.440 152.145 296.570 153.240 ;
        RECT 4.845 147.715 5.975 148.430 ;
        RECT 4.845 147.015 6.000 147.715 ;
        RECT 295.440 147.460 296.570 148.515 ;
        RECT 295.300 147.180 296.570 147.460 ;
        RECT 4.845 146.000 5.975 147.015 ;
        RECT 295.440 146.085 296.570 147.180 ;
        RECT 4.845 141.655 5.975 142.370 ;
        RECT 4.845 140.955 6.000 141.655 ;
        RECT 295.440 141.400 296.570 142.455 ;
        RECT 295.300 141.120 296.570 141.400 ;
        RECT 4.845 139.940 5.975 140.955 ;
        RECT 295.440 140.025 296.570 141.120 ;
        RECT 4.845 135.595 5.975 136.310 ;
        RECT 4.845 134.895 6.000 135.595 ;
        RECT 295.440 135.340 296.570 136.395 ;
        RECT 295.300 135.060 296.570 135.340 ;
        RECT 4.845 133.880 5.975 134.895 ;
        RECT 295.440 133.965 296.570 135.060 ;
        RECT 4.845 129.535 5.975 130.250 ;
        RECT 4.845 128.835 6.000 129.535 ;
        RECT 295.440 129.280 296.570 130.335 ;
        RECT 295.300 129.000 296.570 129.280 ;
        RECT 4.845 127.820 5.975 128.835 ;
        RECT 295.440 127.905 296.570 129.000 ;
        RECT 4.845 123.475 5.975 124.190 ;
        RECT 4.845 122.775 6.000 123.475 ;
        RECT 295.440 123.220 296.570 124.275 ;
        RECT 295.300 122.940 296.570 123.220 ;
        RECT 4.845 121.760 5.975 122.775 ;
        RECT 295.440 121.845 296.570 122.940 ;
        RECT 4.845 117.415 5.975 118.130 ;
        RECT 4.845 116.715 6.000 117.415 ;
        RECT 295.440 117.160 296.570 118.215 ;
        RECT 295.300 116.880 296.570 117.160 ;
        RECT 4.845 115.700 5.975 116.715 ;
        RECT 295.440 115.785 296.570 116.880 ;
        RECT 93.700 5.990 95.245 6.000 ;
      LAYER Metal2 ;
        RECT 2.470 318.940 298.830 319.090 ;
        RECT 2.465 315.890 298.830 318.940 ;
        RECT 2.465 315.590 6.000 315.890 ;
        RECT 295.300 315.590 298.830 315.890 ;
        RECT 2.465 312.050 5.970 315.590 ;
        RECT 295.445 312.270 298.830 315.590 ;
        RECT 2.465 309.620 5.975 312.050 ;
        RECT 2.465 305.990 5.970 309.620 ;
        RECT 2.465 303.560 5.975 305.990 ;
        RECT 2.465 299.930 5.970 303.560 ;
        RECT 2.465 297.500 5.975 299.930 ;
        RECT 2.465 293.870 5.970 297.500 ;
        RECT 2.465 291.440 5.975 293.870 ;
        RECT 2.465 287.810 5.970 291.440 ;
        RECT 2.465 285.380 5.975 287.810 ;
        RECT 2.465 281.750 5.970 285.380 ;
        RECT 2.465 279.320 5.975 281.750 ;
        RECT 2.465 275.690 5.970 279.320 ;
        RECT 2.465 273.260 5.975 275.690 ;
        RECT 2.465 269.630 5.970 273.260 ;
        RECT 2.465 267.200 5.975 269.630 ;
        RECT 2.465 263.570 5.970 267.200 ;
        RECT 2.465 261.140 5.975 263.570 ;
        RECT 2.465 257.510 5.970 261.140 ;
        RECT 2.465 255.080 5.975 257.510 ;
        RECT 2.465 251.450 5.970 255.080 ;
        RECT 2.465 249.020 5.975 251.450 ;
        RECT 2.465 245.390 5.970 249.020 ;
        RECT 2.465 242.960 5.975 245.390 ;
        RECT 2.465 239.330 5.970 242.960 ;
        RECT 2.465 236.900 5.975 239.330 ;
        RECT 2.465 233.270 5.970 236.900 ;
        RECT 2.465 230.840 5.975 233.270 ;
        RECT 2.465 227.210 5.970 230.840 ;
        RECT 2.465 224.780 5.975 227.210 ;
        RECT 2.465 221.150 5.970 224.780 ;
        RECT 2.465 218.720 5.975 221.150 ;
        RECT 2.465 215.090 5.970 218.720 ;
        RECT 2.465 212.660 5.975 215.090 ;
        RECT 2.465 209.030 5.970 212.660 ;
        RECT 2.465 206.600 5.975 209.030 ;
        RECT 2.465 202.970 5.970 206.600 ;
        RECT 2.465 200.540 5.975 202.970 ;
        RECT 2.465 196.910 5.970 200.540 ;
        RECT 2.465 194.480 5.975 196.910 ;
        RECT 2.465 190.850 5.970 194.480 ;
        RECT 2.465 188.420 5.975 190.850 ;
        RECT 2.465 184.790 5.970 188.420 ;
        RECT 2.465 182.360 5.975 184.790 ;
        RECT 2.465 178.730 5.970 182.360 ;
        RECT 2.465 176.300 5.975 178.730 ;
        RECT 2.465 172.670 5.970 176.300 ;
        RECT 2.465 170.240 5.975 172.670 ;
        RECT 2.465 166.610 5.970 170.240 ;
        RECT 295.440 168.360 298.830 312.270 ;
        RECT 2.465 164.180 5.975 166.610 ;
        RECT 2.465 160.550 5.970 164.180 ;
        RECT 2.465 158.120 5.975 160.550 ;
        RECT 2.465 154.490 5.970 158.120 ;
        RECT 2.465 152.060 5.975 154.490 ;
        RECT 2.465 148.430 5.970 152.060 ;
        RECT 2.465 146.000 5.975 148.430 ;
        RECT 2.465 142.370 5.970 146.000 ;
        RECT 2.465 139.940 5.975 142.370 ;
        RECT 2.465 136.310 5.970 139.940 ;
        RECT 2.465 133.880 5.975 136.310 ;
        RECT 2.465 130.250 5.970 133.880 ;
        RECT 2.465 127.820 5.975 130.250 ;
        RECT 2.465 124.190 5.970 127.820 ;
        RECT 2.465 121.760 5.975 124.190 ;
        RECT 2.465 118.130 5.970 121.760 ;
        RECT 2.465 115.700 5.975 118.130 ;
        RECT 2.465 110.435 5.970 115.700 ;
        RECT 295.440 110.435 298.835 168.360 ;
        RECT 2.465 4.330 5.975 110.435 ;
        RECT 26.795 4.830 27.580 6.000 ;
        RECT 65.605 4.830 66.390 6.000 ;
        RECT 2.465 1.410 5.970 4.330 ;
        RECT 88.750 4.285 89.535 6.000 ;
        RECT 93.695 5.965 95.245 6.000 ;
        RECT 131.250 5.180 132.035 6.000 ;
        RECT 137.620 5.180 138.405 6.000 ;
        RECT 207.850 4.315 208.635 6.000 ;
        RECT 232.070 4.830 232.855 6.000 ;
        RECT 271.220 4.810 272.005 6.000 ;
        RECT 295.330 4.330 298.835 110.435 ;
        RECT 2.470 0.985 5.970 1.410 ;
        RECT 295.330 0.985 298.830 4.330 ;
      LAYER Metal3 ;
        RECT 5.090 319.760 8.590 321.890 ;
        RECT 5.090 319.090 8.585 319.760 ;
        RECT 14.480 319.090 17.975 321.890 ;
        RECT 24.630 319.760 28.130 321.890 ;
        RECT 33.380 321.190 36.880 321.890 ;
        RECT 24.630 319.090 28.125 319.760 ;
        RECT 33.380 319.090 36.875 321.190 ;
        RECT 44.170 319.090 47.665 321.890 ;
        RECT 52.280 319.090 55.775 321.890 ;
        RECT 63.710 319.090 67.205 321.890 ;
        RECT 72.285 319.090 75.780 321.890 ;
        RECT 84.680 319.760 88.180 321.890 ;
        RECT 84.685 319.090 88.180 319.760 ;
        RECT 93.000 319.090 96.495 321.890 ;
        RECT 107.485 319.090 110.980 321.890 ;
        RECT 123.950 319.090 127.445 321.890 ;
        RECT 135.045 319.090 138.540 321.890 ;
        RECT 144.305 319.090 147.800 321.890 ;
        RECT 157.740 319.090 161.235 321.890 ;
        RECT 162.095 319.090 165.590 321.890 ;
        RECT 171.155 319.090 174.650 321.890 ;
        RECT 183.990 319.090 187.485 321.890 ;
        RECT 189.915 319.090 193.410 321.890 ;
        RECT 201.415 319.090 204.910 321.890 ;
        RECT 210.520 319.090 214.015 321.890 ;
        RECT 221.995 319.090 225.490 321.890 ;
        RECT 230.060 319.090 233.555 321.890 ;
        RECT 240.895 319.090 244.390 321.890 ;
        RECT 249.600 319.090 253.095 321.890 ;
        RECT 259.795 319.090 263.290 321.890 ;
        RECT 269.125 319.090 272.620 321.890 ;
        RECT 279.300 319.090 282.795 321.890 ;
        RECT 290.115 319.090 293.610 321.890 ;
        RECT 295.330 319.090 298.825 321.890 ;
        RECT 0.000 315.890 301.300 319.090 ;
        RECT 0.000 315.590 6.000 315.890 ;
        RECT 295.300 315.590 301.300 315.890 ;
        RECT 5.090 315.585 6.000 315.590 ;
        RECT 296.440 312.135 301.300 312.145 ;
        RECT 0.000 309.610 5.975 312.060 ;
        RECT 295.440 309.705 301.300 312.135 ;
        RECT 296.440 309.695 301.300 309.705 ;
        RECT 296.440 306.075 301.300 306.085 ;
        RECT 0.000 303.550 5.975 306.000 ;
        RECT 295.440 303.645 301.300 306.075 ;
        RECT 296.440 303.635 301.300 303.645 ;
        RECT 296.440 300.015 301.300 300.025 ;
        RECT 0.000 297.490 5.975 299.940 ;
        RECT 295.440 297.585 301.300 300.015 ;
        RECT 296.440 297.575 301.300 297.585 ;
        RECT 296.440 293.955 301.300 293.965 ;
        RECT 0.000 291.430 5.975 293.880 ;
        RECT 295.440 291.525 301.300 293.955 ;
        RECT 296.440 291.515 301.300 291.525 ;
        RECT 296.440 287.895 301.300 287.905 ;
        RECT 0.000 285.370 5.975 287.820 ;
        RECT 295.440 285.465 301.300 287.895 ;
        RECT 296.440 285.455 301.300 285.465 ;
        RECT 296.440 281.835 301.300 281.845 ;
        RECT 0.000 279.310 5.975 281.760 ;
        RECT 295.440 279.405 301.300 281.835 ;
        RECT 296.440 279.395 301.300 279.405 ;
        RECT 296.440 275.775 301.300 275.785 ;
        RECT 0.000 273.250 5.975 275.700 ;
        RECT 295.440 273.345 301.300 275.775 ;
        RECT 296.440 273.335 301.300 273.345 ;
        RECT 296.440 269.715 301.300 269.725 ;
        RECT 0.000 267.190 5.975 269.640 ;
        RECT 295.440 267.285 301.300 269.715 ;
        RECT 296.440 267.275 301.300 267.285 ;
        RECT 296.440 263.655 301.300 263.665 ;
        RECT 0.000 261.130 5.975 263.580 ;
        RECT 295.440 261.225 301.300 263.655 ;
        RECT 296.440 261.215 301.300 261.225 ;
        RECT 296.440 257.595 301.300 257.605 ;
        RECT 0.000 255.070 5.975 257.520 ;
        RECT 295.440 255.165 301.300 257.595 ;
        RECT 296.440 255.155 301.300 255.165 ;
        RECT 296.440 251.535 301.300 251.545 ;
        RECT 0.000 249.010 5.975 251.460 ;
        RECT 295.440 249.105 301.300 251.535 ;
        RECT 296.440 249.095 301.300 249.105 ;
        RECT 296.440 245.475 301.300 245.485 ;
        RECT 0.000 242.950 5.975 245.400 ;
        RECT 295.440 243.045 301.300 245.475 ;
        RECT 296.440 243.035 301.300 243.045 ;
        RECT 296.440 239.415 301.300 239.425 ;
        RECT 0.000 236.890 5.975 239.340 ;
        RECT 295.440 236.985 301.300 239.415 ;
        RECT 296.440 236.975 301.300 236.985 ;
        RECT 296.440 233.355 301.300 233.365 ;
        RECT 0.000 230.830 5.975 233.280 ;
        RECT 295.440 230.925 301.300 233.355 ;
        RECT 296.440 230.915 301.300 230.925 ;
        RECT 296.440 227.295 301.300 227.305 ;
        RECT 0.000 224.770 5.975 227.220 ;
        RECT 295.440 224.865 301.300 227.295 ;
        RECT 296.440 224.855 301.300 224.865 ;
        RECT 296.440 221.235 301.300 221.245 ;
        RECT 0.000 218.710 5.975 221.160 ;
        RECT 295.440 218.805 301.300 221.235 ;
        RECT 296.440 218.795 301.300 218.805 ;
        RECT 296.440 215.175 301.300 215.185 ;
        RECT 0.000 212.650 5.975 215.100 ;
        RECT 295.440 212.745 301.300 215.175 ;
        RECT 296.440 212.735 301.300 212.745 ;
        RECT 296.440 209.115 301.300 209.125 ;
        RECT 0.000 206.590 5.975 209.040 ;
        RECT 295.440 206.685 301.300 209.115 ;
        RECT 296.440 206.675 301.300 206.685 ;
        RECT 296.440 203.055 301.300 203.065 ;
        RECT 0.000 200.530 5.975 202.980 ;
        RECT 295.440 200.625 301.300 203.055 ;
        RECT 296.440 200.615 301.300 200.625 ;
        RECT 296.440 196.995 301.300 197.005 ;
        RECT 0.000 194.470 5.975 196.920 ;
        RECT 295.440 194.565 301.300 196.995 ;
        RECT 296.440 194.555 301.300 194.565 ;
        RECT 296.440 190.935 301.300 190.945 ;
        RECT 0.000 188.410 5.975 190.860 ;
        RECT 295.440 188.505 301.300 190.935 ;
        RECT 296.440 188.495 301.300 188.505 ;
        RECT 296.440 184.875 301.300 184.885 ;
        RECT 0.000 182.350 5.975 184.800 ;
        RECT 295.440 182.445 301.300 184.875 ;
        RECT 296.440 182.435 301.300 182.445 ;
        RECT 296.440 178.815 301.300 178.825 ;
        RECT 0.000 176.290 5.975 178.740 ;
        RECT 295.440 176.385 301.300 178.815 ;
        RECT 296.440 176.375 301.300 176.385 ;
        RECT 296.440 172.755 301.300 172.765 ;
        RECT 0.000 170.230 5.975 172.680 ;
        RECT 295.440 170.325 301.300 172.755 ;
        RECT 296.440 170.315 301.300 170.325 ;
        RECT 296.440 166.695 301.300 166.705 ;
        RECT 0.000 164.170 5.975 166.620 ;
        RECT 295.440 164.265 301.300 166.695 ;
        RECT 296.440 164.255 301.300 164.265 ;
        RECT 296.440 160.635 301.300 160.645 ;
        RECT 0.000 158.110 5.975 160.560 ;
        RECT 295.440 158.205 301.300 160.635 ;
        RECT 296.440 158.195 301.300 158.205 ;
        RECT 296.440 154.575 301.300 154.585 ;
        RECT 0.000 152.050 5.975 154.500 ;
        RECT 295.440 152.145 301.300 154.575 ;
        RECT 296.440 152.135 301.300 152.145 ;
        RECT 296.440 148.515 301.300 148.525 ;
        RECT 0.000 145.990 5.975 148.440 ;
        RECT 295.440 146.085 301.300 148.515 ;
        RECT 296.440 146.075 301.300 146.085 ;
        RECT 296.440 142.455 301.300 142.465 ;
        RECT 0.000 139.930 5.975 142.380 ;
        RECT 295.440 140.025 301.300 142.455 ;
        RECT 296.440 140.015 301.300 140.025 ;
        RECT 296.440 136.395 301.300 136.405 ;
        RECT 0.000 133.870 5.975 136.320 ;
        RECT 295.440 133.965 301.300 136.395 ;
        RECT 296.440 133.955 301.300 133.965 ;
        RECT 296.440 130.335 301.300 130.345 ;
        RECT 0.000 127.810 5.975 130.260 ;
        RECT 295.440 127.905 301.300 130.335 ;
        RECT 296.440 127.895 301.300 127.905 ;
        RECT 296.440 124.275 301.300 124.285 ;
        RECT 0.000 121.750 5.975 124.200 ;
        RECT 295.440 121.845 301.300 124.275 ;
        RECT 296.440 121.835 301.300 121.845 ;
        RECT 296.440 118.215 301.300 118.225 ;
        RECT 0.000 115.690 5.975 118.140 ;
        RECT 295.440 115.785 301.300 118.215 ;
        RECT 296.440 115.775 301.300 115.785 ;
        RECT 0.000 109.905 3.545 109.910 ;
        RECT 297.750 109.905 301.300 109.910 ;
        RECT 0.000 102.880 6.000 109.905 ;
        RECT 295.300 102.880 301.300 109.905 ;
        RECT 0.000 96.170 5.975 102.880 ;
        RECT 295.335 96.170 301.300 102.880 ;
        RECT 0.000 95.175 6.000 96.170 ;
        RECT 295.300 95.175 301.300 96.170 ;
        RECT 300.600 95.170 301.300 95.175 ;
        RECT 0.000 78.350 3.545 78.355 ;
        RECT 297.750 78.350 301.300 78.355 ;
        RECT 0.000 76.400 5.975 78.350 ;
        RECT 295.335 76.400 301.300 78.350 ;
        RECT 0.000 74.855 6.000 76.400 ;
        RECT 0.010 74.850 6.000 74.855 ;
        RECT 295.300 74.850 301.300 76.400 ;
        RECT 297.750 67.740 301.300 67.750 ;
        RECT 0.010 67.735 6.000 67.740 ;
        RECT 0.000 58.210 6.000 67.735 ;
        RECT 295.300 58.210 301.300 67.740 ;
        RECT 0.000 58.205 0.700 58.210 ;
        RECT 300.600 58.205 301.300 58.210 ;
        RECT 0.000 47.315 3.545 47.325 ;
        RECT 300.600 47.315 301.300 47.320 ;
        RECT 0.000 44.810 6.000 47.315 ;
        RECT 295.300 44.810 301.300 47.315 ;
        RECT 0.000 42.955 5.975 44.810 ;
        RECT 295.335 42.970 301.300 44.810 ;
        RECT 0.000 40.125 6.000 42.955 ;
        RECT 0.010 40.120 6.000 40.125 ;
        RECT 295.300 40.120 301.300 42.970 ;
        RECT 0.010 40.020 5.975 40.120 ;
        RECT 295.335 40.020 301.300 40.120 ;
        RECT 297.750 40.010 301.300 40.020 ;
        RECT 0.000 31.295 3.545 31.300 ;
        RECT 295.300 31.295 295.365 31.325 ;
        RECT 300.600 31.295 301.300 31.300 ;
        RECT 0.000 26.530 6.000 31.295 ;
        RECT 0.010 26.525 6.000 26.530 ;
        RECT 295.300 26.525 301.300 31.295 ;
        RECT 0.000 19.345 3.545 19.350 ;
        RECT 297.750 19.345 301.300 19.350 ;
        RECT 0.000 17.750 6.000 19.345 ;
        RECT 0.000 15.795 5.995 17.750 ;
        RECT 295.300 17.745 301.300 19.345 ;
        RECT 295.315 15.805 301.300 17.745 ;
        RECT 0.000 14.210 6.000 15.795 ;
        RECT 0.010 14.205 6.000 14.210 ;
        RECT 295.300 14.205 301.300 15.805 ;
        RECT 0.000 6.000 6.000 7.810 ;
        RECT 295.300 6.000 301.300 7.810 ;
        RECT 0.000 4.310 301.300 6.000 ;
        RECT 0.000 4.290 0.700 4.310 ;
        RECT 2.465 0.000 5.970 4.310 ;
        RECT 7.135 0.000 10.635 4.310 ;
        RECT 12.045 0.000 15.545 4.310 ;
        RECT 20.445 0.000 23.945 4.310 ;
        RECT 24.645 0.000 28.145 4.310 ;
        RECT 28.845 0.000 32.345 4.310 ;
        RECT 37.245 0.000 40.745 4.310 ;
        RECT 43.550 0.000 47.050 4.310 ;
        RECT 49.845 0.000 53.345 4.310 ;
        RECT 58.245 0.000 61.745 4.310 ;
        RECT 62.445 0.000 65.945 4.310 ;
        RECT 66.645 0.000 70.145 4.310 ;
        RECT 76.685 0.000 80.185 4.310 ;
        RECT 80.885 0.000 84.385 4.310 ;
        RECT 85.435 0.000 88.935 4.310 ;
        RECT 89.985 0.000 93.485 4.310 ;
        RECT 94.535 0.000 98.035 4.310 ;
        RECT 99.085 0.000 102.585 4.310 ;
        RECT 103.635 0.000 107.135 4.310 ;
        RECT 126.105 0.000 129.605 4.310 ;
        RECT 137.295 0.000 140.795 4.310 ;
        RECT 148.515 0.000 152.015 4.310 ;
        RECT 156.915 0.000 160.415 4.310 ;
        RECT 165.315 0.000 168.815 4.310 ;
        RECT 169.980 0.000 173.480 4.310 ;
        RECT 174.565 0.000 178.065 4.310 ;
        RECT 190.600 0.000 194.100 4.310 ;
        RECT 195.150 0.000 198.650 4.310 ;
        RECT 199.700 4.205 221.530 4.310 ;
        RECT 199.700 0.000 203.200 4.205 ;
        RECT 204.250 0.000 207.750 4.205 ;
        RECT 208.800 0.000 212.300 4.205 ;
        RECT 213.350 0.000 216.850 4.205 ;
        RECT 218.030 0.000 221.530 4.205 ;
        RECT 227.960 0.000 231.460 4.310 ;
        RECT 232.160 0.000 235.660 4.310 ;
        RECT 236.360 0.000 239.860 4.310 ;
        RECT 244.760 0.000 248.260 4.310 ;
        RECT 251.055 0.000 254.555 4.310 ;
        RECT 257.360 0.000 260.860 4.310 ;
        RECT 265.760 0.000 269.260 4.310 ;
        RECT 269.960 0.000 273.460 4.310 ;
        RECT 274.160 0.000 277.660 4.310 ;
        RECT 283.560 0.000 287.060 4.310 ;
        RECT 288.465 0.000 291.965 4.310 ;
        RECT 295.330 0.000 298.830 4.310 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.985 317.365 300.315 320.900 ;
        RECT 0.985 315.035 4.485 317.365 ;
        RECT 7.150 315.890 7.970 317.365 ;
        RECT 26.690 315.890 27.510 317.365 ;
        RECT 46.230 315.890 47.050 317.365 ;
        RECT 65.770 315.890 66.590 317.365 ;
        RECT 85.300 315.890 86.120 317.365 ;
        RECT 90.140 315.890 92.685 317.365 ;
        RECT 96.620 317.030 102.185 317.365 ;
        RECT 95.855 315.890 102.185 317.030 ;
        RECT 119.790 315.890 122.545 317.365 ;
        RECT 140.215 315.890 142.065 317.365 ;
        RECT 153.080 315.890 155.970 317.365 ;
        RECT 175.340 315.890 178.195 317.365 ;
        RECT 194.845 315.890 202.075 317.365 ;
        RECT 204.765 315.890 207.310 317.365 ;
        RECT 212.580 315.890 213.400 317.365 ;
        RECT 232.120 315.890 232.940 317.365 ;
        RECT 251.660 315.890 252.480 317.365 ;
        RECT 271.185 315.890 272.005 317.365 ;
        RECT 290.730 315.890 291.550 317.365 ;
        RECT 0.985 314.885 4.490 315.035 ;
        RECT 0.985 313.080 6.000 314.885 ;
        RECT 0.985 309.785 4.490 313.080 ;
        RECT 0.985 308.975 4.485 309.785 ;
        RECT 0.985 308.825 4.490 308.975 ;
        RECT 0.985 307.020 6.000 308.825 ;
        RECT 0.985 303.725 4.490 307.020 ;
        RECT 0.985 302.915 4.485 303.725 ;
        RECT 0.985 302.765 4.490 302.915 ;
        RECT 0.985 300.960 6.000 302.765 ;
        RECT 0.985 297.665 4.490 300.960 ;
        RECT 0.985 296.855 4.485 297.665 ;
        RECT 0.985 296.705 4.490 296.855 ;
        RECT 0.985 294.900 6.000 296.705 ;
        RECT 0.985 291.605 4.490 294.900 ;
        RECT 0.985 290.795 4.485 291.605 ;
        RECT 0.985 290.645 4.490 290.795 ;
        RECT 0.985 288.840 6.000 290.645 ;
        RECT 295.300 289.410 296.325 290.110 ;
        RECT 0.985 285.545 4.490 288.840 ;
        RECT 0.985 284.735 4.485 285.545 ;
        RECT 0.985 284.585 4.490 284.735 ;
        RECT 0.985 282.780 6.000 284.585 ;
        RECT 0.985 279.485 4.490 282.780 ;
        RECT 0.985 278.675 4.485 279.485 ;
        RECT 0.985 278.525 4.490 278.675 ;
        RECT 0.985 276.720 6.000 278.525 ;
        RECT 0.985 273.425 4.490 276.720 ;
        RECT 0.985 272.615 4.485 273.425 ;
        RECT 0.985 272.465 4.490 272.615 ;
        RECT 0.985 270.660 6.000 272.465 ;
        RECT 0.985 267.365 4.490 270.660 ;
        RECT 0.985 266.555 4.485 267.365 ;
        RECT 0.985 266.405 4.490 266.555 ;
        RECT 0.985 264.600 6.000 266.405 ;
        RECT 0.985 261.305 4.490 264.600 ;
        RECT 0.985 260.495 4.485 261.305 ;
        RECT 0.985 260.345 4.490 260.495 ;
        RECT 0.985 258.540 6.000 260.345 ;
        RECT 0.985 255.245 4.490 258.540 ;
        RECT 0.985 254.435 4.485 255.245 ;
        RECT 0.985 254.285 4.490 254.435 ;
        RECT 0.985 252.480 6.000 254.285 ;
        RECT 0.985 249.185 4.490 252.480 ;
        RECT 0.985 248.375 4.485 249.185 ;
        RECT 0.985 248.225 4.490 248.375 ;
        RECT 0.985 246.420 6.000 248.225 ;
        RECT 0.985 243.125 4.490 246.420 ;
        RECT 0.985 242.315 4.485 243.125 ;
        RECT 0.985 242.165 4.490 242.315 ;
        RECT 0.985 240.360 6.000 242.165 ;
        RECT 0.985 237.065 4.490 240.360 ;
        RECT 0.985 236.255 4.485 237.065 ;
        RECT 0.985 236.105 4.490 236.255 ;
        RECT 0.985 234.300 6.000 236.105 ;
        RECT 0.985 231.005 4.490 234.300 ;
        RECT 0.985 230.195 4.485 231.005 ;
        RECT 0.985 230.045 4.490 230.195 ;
        RECT 0.985 228.240 6.000 230.045 ;
        RECT 0.985 224.945 4.490 228.240 ;
        RECT 0.985 224.135 4.485 224.945 ;
        RECT 0.985 223.985 4.490 224.135 ;
        RECT 0.985 222.180 6.000 223.985 ;
        RECT 0.985 218.885 4.490 222.180 ;
        RECT 0.985 218.075 4.485 218.885 ;
        RECT 0.985 217.925 4.490 218.075 ;
        RECT 0.985 216.120 6.000 217.925 ;
        RECT 0.985 212.825 4.490 216.120 ;
        RECT 0.985 212.015 4.485 212.825 ;
        RECT 0.985 211.865 4.490 212.015 ;
        RECT 0.985 210.060 6.000 211.865 ;
        RECT 0.985 206.765 4.490 210.060 ;
        RECT 0.985 205.955 4.485 206.765 ;
        RECT 0.985 205.805 4.490 205.955 ;
        RECT 0.985 204.000 6.000 205.805 ;
        RECT 0.985 200.705 4.490 204.000 ;
        RECT 0.985 199.895 4.485 200.705 ;
        RECT 0.985 199.745 4.490 199.895 ;
        RECT 0.985 197.940 6.000 199.745 ;
        RECT 0.985 194.645 4.490 197.940 ;
        RECT 0.985 193.835 4.485 194.645 ;
        RECT 0.985 193.685 4.490 193.835 ;
        RECT 0.985 191.880 6.000 193.685 ;
        RECT 0.985 188.585 4.490 191.880 ;
        RECT 0.985 187.775 4.485 188.585 ;
        RECT 0.985 187.625 4.490 187.775 ;
        RECT 0.985 185.820 6.000 187.625 ;
        RECT 0.985 182.525 4.490 185.820 ;
        RECT 0.985 181.715 4.485 182.525 ;
        RECT 0.985 181.565 4.490 181.715 ;
        RECT 0.985 179.760 6.000 181.565 ;
        RECT 0.985 176.465 4.490 179.760 ;
        RECT 0.985 175.655 4.485 176.465 ;
        RECT 0.985 175.505 4.490 175.655 ;
        RECT 0.985 173.700 6.000 175.505 ;
        RECT 0.985 170.405 4.490 173.700 ;
        RECT 0.985 169.595 4.485 170.405 ;
        RECT 0.985 169.445 4.490 169.595 ;
        RECT 0.985 167.640 6.000 169.445 ;
        RECT 0.985 164.345 4.490 167.640 ;
        RECT 0.985 163.535 4.485 164.345 ;
        RECT 0.985 163.385 4.490 163.535 ;
        RECT 0.985 161.580 6.000 163.385 ;
        RECT 0.985 158.285 4.490 161.580 ;
        RECT 0.985 157.475 4.485 158.285 ;
        RECT 0.985 157.325 4.490 157.475 ;
        RECT 0.985 155.520 6.000 157.325 ;
        RECT 0.985 152.225 4.490 155.520 ;
        RECT 0.985 151.415 4.485 152.225 ;
        RECT 0.985 151.265 4.490 151.415 ;
        RECT 0.985 149.460 6.000 151.265 ;
        RECT 0.985 146.165 4.490 149.460 ;
        RECT 0.985 145.355 4.485 146.165 ;
        RECT 0.985 145.205 4.490 145.355 ;
        RECT 0.985 143.400 6.000 145.205 ;
        RECT 0.985 140.105 4.490 143.400 ;
        RECT 0.985 139.295 4.485 140.105 ;
        RECT 0.985 139.145 4.490 139.295 ;
        RECT 0.985 137.340 6.000 139.145 ;
        RECT 0.985 134.045 4.490 137.340 ;
        RECT 0.985 133.235 4.485 134.045 ;
        RECT 0.985 133.085 4.490 133.235 ;
        RECT 0.985 131.280 6.000 133.085 ;
        RECT 0.985 127.985 4.490 131.280 ;
        RECT 0.985 127.175 4.485 127.985 ;
        RECT 0.985 127.025 4.490 127.175 ;
        RECT 0.985 125.220 6.000 127.025 ;
        RECT 0.985 121.925 4.490 125.220 ;
        RECT 0.985 121.115 4.485 121.925 ;
        RECT 0.985 120.965 4.490 121.115 ;
        RECT 0.985 119.160 6.000 120.965 ;
        RECT 0.985 115.865 4.490 119.160 ;
        RECT 0.985 87.265 4.485 115.865 ;
        RECT 296.815 114.965 300.315 317.365 ;
        RECT 295.300 114.355 300.315 114.965 ;
        RECT 296.815 112.405 300.315 114.355 ;
        RECT 295.300 111.810 300.315 112.405 ;
        RECT 296.815 87.265 300.315 111.810 ;
        RECT 0.985 86.795 6.000 87.265 ;
        RECT 295.300 86.795 300.315 87.265 ;
        RECT 0.985 72.515 4.485 86.795 ;
        RECT 296.815 72.515 300.315 86.795 ;
        RECT 0.985 71.835 6.000 72.515 ;
        RECT 295.300 71.835 300.315 72.515 ;
        RECT 0.985 4.485 4.485 71.835 ;
        RECT 95.850 4.485 202.075 6.000 ;
        RECT 296.815 4.485 300.315 71.835 ;
        RECT 0.985 4.480 202.505 4.485 ;
        RECT 204.680 4.480 300.315 4.485 ;
        RECT 0.985 0.985 300.315 4.480 ;
        RECT 87.030 0.980 87.730 0.985 ;
        RECT 90.590 0.980 91.290 0.985 ;
      LAYER Metal2 ;
        RECT 0.985 319.760 300.315 320.900 ;
        RECT 0.995 312.770 2.125 315.200 ;
        RECT 299.120 312.755 300.800 315.185 ;
        RECT 0.995 306.710 2.125 309.140 ;
        RECT 299.120 306.695 300.800 309.125 ;
        RECT 0.995 300.650 2.125 303.080 ;
        RECT 299.120 300.635 300.800 303.065 ;
        RECT 0.995 294.590 2.125 297.020 ;
        RECT 299.120 294.575 300.800 297.005 ;
        RECT 0.995 288.530 2.125 290.960 ;
        RECT 299.120 288.515 300.800 290.945 ;
        RECT 0.995 282.470 2.125 284.900 ;
        RECT 299.120 282.455 300.800 284.885 ;
        RECT 0.995 276.410 2.125 278.840 ;
        RECT 299.120 276.395 300.800 278.825 ;
        RECT 0.995 270.350 2.125 272.780 ;
        RECT 299.120 270.335 300.800 272.765 ;
        RECT 0.995 264.290 2.125 266.720 ;
        RECT 299.120 264.275 300.800 266.705 ;
        RECT 0.995 258.230 2.125 260.660 ;
        RECT 299.120 258.215 300.800 260.645 ;
        RECT 0.995 252.170 2.125 254.600 ;
        RECT 299.120 252.155 300.800 254.585 ;
        RECT 0.995 246.110 2.125 248.540 ;
        RECT 299.120 246.095 300.800 248.525 ;
        RECT 0.995 240.050 2.125 242.480 ;
        RECT 299.120 240.035 300.800 242.465 ;
        RECT 0.995 233.990 2.125 236.420 ;
        RECT 299.120 233.975 300.800 236.405 ;
        RECT 0.995 227.930 2.125 230.360 ;
        RECT 299.120 227.915 300.800 230.345 ;
        RECT 0.995 221.870 2.125 224.300 ;
        RECT 299.120 221.855 300.800 224.285 ;
        RECT 0.995 215.810 2.125 218.240 ;
        RECT 299.120 215.795 300.800 218.225 ;
        RECT 0.995 209.750 2.125 212.180 ;
        RECT 299.120 209.735 300.800 212.165 ;
        RECT 0.995 203.690 2.125 206.120 ;
        RECT 299.120 203.675 300.800 206.105 ;
        RECT 0.995 197.630 2.125 200.060 ;
        RECT 299.120 197.615 300.800 200.045 ;
        RECT 0.995 191.570 2.125 194.000 ;
        RECT 299.120 191.555 300.800 193.985 ;
        RECT 0.995 185.510 2.125 187.940 ;
        RECT 299.120 185.495 300.800 187.925 ;
        RECT 0.995 179.450 2.125 181.880 ;
        RECT 299.120 179.435 300.800 181.865 ;
        RECT 0.995 173.390 2.125 175.820 ;
        RECT 299.120 173.375 300.800 175.805 ;
        RECT 0.995 167.330 2.125 169.760 ;
        RECT 299.120 167.315 300.800 169.745 ;
        RECT 0.995 161.270 2.125 163.700 ;
        RECT 299.120 161.255 300.800 163.685 ;
        RECT 0.995 155.210 2.125 157.640 ;
        RECT 299.120 155.195 300.800 157.625 ;
        RECT 0.995 149.150 2.125 151.580 ;
        RECT 299.120 149.135 300.800 151.565 ;
        RECT 0.995 143.090 2.125 145.520 ;
        RECT 299.120 143.075 300.800 145.505 ;
        RECT 0.995 137.030 2.125 139.460 ;
        RECT 299.120 137.015 300.800 139.445 ;
        RECT 0.995 130.970 2.125 133.400 ;
        RECT 299.120 130.955 300.800 133.385 ;
        RECT 0.995 124.910 2.125 127.340 ;
        RECT 299.120 124.895 300.800 127.325 ;
        RECT 0.995 118.850 2.125 121.280 ;
        RECT 299.120 118.835 300.800 121.265 ;
        RECT 0.995 111.495 2.125 113.925 ;
        RECT 299.185 111.495 300.315 113.925 ;
        RECT 0.995 83.455 2.125 92.695 ;
        RECT 299.185 83.455 300.315 92.695 ;
        RECT 0.995 69.460 2.125 72.760 ;
        RECT 299.185 69.460 300.315 72.760 ;
        RECT 0.995 48.095 2.125 57.145 ;
        RECT 299.185 48.095 300.315 57.145 ;
        RECT 0.995 33.790 2.125 37.960 ;
        RECT 299.185 33.790 300.315 37.960 ;
        RECT 0.995 19.880 2.125 26.220 ;
        RECT 299.185 19.880 300.315 26.220 ;
        RECT 0.995 8.890 2.125 13.060 ;
        RECT 299.185 8.890 300.315 13.060 ;
        RECT 16.245 0.985 19.745 4.485 ;
        RECT 25.040 0.985 25.820 6.000 ;
        RECT 28.600 0.985 29.385 6.000 ;
        RECT 33.045 0.985 36.545 4.485 ;
        RECT 54.045 0.985 57.545 4.485 ;
        RECT 63.850 0.985 64.630 6.000 ;
        RECT 67.410 0.985 68.195 6.000 ;
        RECT 70.845 0.985 74.345 4.485 ;
        RECT 87.000 0.975 87.775 6.000 ;
        RECT 90.555 0.975 91.335 6.000 ;
        RECT 109.630 0.985 113.130 4.485 ;
        RECT 115.575 0.985 119.075 4.485 ;
        RECT 121.905 0.985 125.405 4.485 ;
        RECT 129.495 4.310 130.275 6.000 ;
        RECT 133.055 4.485 133.840 6.000 ;
        RECT 135.865 4.485 136.645 6.000 ;
        RECT 133.055 4.310 136.645 4.485 ;
        RECT 139.425 4.310 140.210 6.000 ;
        RECT 133.095 0.985 136.595 4.310 ;
        RECT 144.315 0.985 147.815 4.485 ;
        RECT 152.715 0.985 156.215 4.485 ;
        RECT 161.115 0.985 164.615 4.485 ;
        RECT 179.315 0.985 182.815 4.485 ;
        RECT 183.670 0.985 187.170 4.485 ;
        RECT 206.100 1.005 206.875 6.000 ;
        RECT 209.655 1.005 210.435 6.000 ;
        RECT 223.760 0.985 227.260 4.485 ;
        RECT 230.315 0.985 231.095 6.000 ;
        RECT 233.875 0.985 234.660 6.000 ;
        RECT 240.560 0.985 244.060 4.485 ;
        RECT 261.560 0.985 265.060 4.485 ;
        RECT 269.465 0.965 270.245 6.000 ;
        RECT 273.025 0.965 273.810 6.000 ;
        RECT 278.360 0.985 281.860 4.485 ;
      LAYER Metal3 ;
        RECT 9.370 319.755 12.870 321.890 ;
        RECT 18.760 319.760 22.260 321.890 ;
        RECT 28.910 319.755 32.410 321.890 ;
        RECT 37.660 319.760 41.160 321.890 ;
        RECT 48.450 319.755 51.950 321.890 ;
        RECT 56.560 319.760 60.060 321.890 ;
        RECT 67.990 319.755 71.490 321.890 ;
        RECT 80.400 319.755 83.900 321.890 ;
        RECT 88.805 319.760 92.305 321.890 ;
        RECT 98.320 319.760 101.820 321.890 ;
        RECT 103.205 319.760 106.705 321.890 ;
        RECT 114.085 319.760 117.585 321.890 ;
        RECT 119.835 319.760 123.335 321.890 ;
        RECT 130.070 319.760 133.570 321.890 ;
        RECT 140.340 319.760 143.840 321.890 ;
        RECT 149.255 319.760 152.755 321.890 ;
        RECT 153.745 319.760 157.245 321.890 ;
        RECT 166.375 319.760 169.875 321.890 ;
        RECT 177.380 319.760 180.880 321.890 ;
        RECT 196.715 319.760 200.215 321.890 ;
        RECT 205.520 319.760 209.020 321.890 ;
        RECT 214.800 319.755 218.300 321.890 ;
        RECT 226.275 319.760 229.775 321.890 ;
        RECT 234.340 319.755 237.840 321.890 ;
        RECT 245.175 319.760 248.675 321.890 ;
        RECT 253.880 319.755 257.380 321.890 ;
        RECT 264.075 319.760 267.575 321.890 ;
        RECT 273.405 319.755 276.905 321.890 ;
        RECT 285.830 319.755 289.330 321.890 ;
        RECT 0.000 314.510 3.555 315.210 ;
        RECT 297.755 315.090 301.300 315.195 ;
        RECT 297.750 314.695 301.300 315.090 ;
        RECT 0.000 313.460 6.000 314.510 ;
        RECT 295.300 313.645 301.300 314.695 ;
        RECT 0.000 312.760 3.555 313.460 ;
        RECT 297.750 312.645 301.300 313.645 ;
        RECT 0.000 308.450 3.555 309.150 ;
        RECT 297.750 308.635 301.300 309.135 ;
        RECT 0.000 307.400 6.000 308.450 ;
        RECT 295.300 307.585 301.300 308.635 ;
        RECT 0.000 306.700 3.555 307.400 ;
        RECT 297.750 306.685 301.300 307.585 ;
        RECT 0.000 302.390 3.555 303.090 ;
        RECT 297.750 302.575 301.300 303.075 ;
        RECT 0.000 301.340 6.000 302.390 ;
        RECT 295.300 301.525 301.300 302.575 ;
        RECT 0.000 300.640 3.555 301.340 ;
        RECT 297.750 300.625 301.300 301.525 ;
        RECT 0.000 296.330 3.555 297.030 ;
        RECT 297.750 296.515 301.300 297.015 ;
        RECT 0.000 295.280 6.000 296.330 ;
        RECT 295.300 295.465 301.300 296.515 ;
        RECT 0.000 294.580 3.555 295.280 ;
        RECT 297.750 294.565 301.300 295.465 ;
        RECT 0.000 290.270 3.555 290.970 ;
        RECT 297.750 290.455 301.300 290.955 ;
        RECT 0.000 289.220 6.000 290.270 ;
        RECT 295.300 289.405 301.300 290.455 ;
        RECT 0.000 288.520 3.555 289.220 ;
        RECT 297.750 288.505 301.300 289.405 ;
        RECT 0.000 284.210 3.555 284.910 ;
        RECT 297.750 284.395 301.300 284.895 ;
        RECT 0.000 283.160 6.000 284.210 ;
        RECT 295.300 283.345 301.300 284.395 ;
        RECT 0.000 282.460 3.555 283.160 ;
        RECT 297.750 282.445 301.300 283.345 ;
        RECT 0.000 278.150 3.555 278.850 ;
        RECT 297.750 278.335 301.300 278.835 ;
        RECT 0.000 277.100 6.000 278.150 ;
        RECT 295.300 277.285 301.300 278.335 ;
        RECT 0.000 276.400 3.555 277.100 ;
        RECT 297.750 276.385 301.300 277.285 ;
        RECT 0.000 272.090 3.555 272.790 ;
        RECT 297.750 272.275 301.300 272.775 ;
        RECT 0.000 271.040 6.000 272.090 ;
        RECT 295.300 271.225 301.300 272.275 ;
        RECT 0.000 270.340 3.555 271.040 ;
        RECT 297.750 270.325 301.300 271.225 ;
        RECT 0.000 266.030 3.555 266.730 ;
        RECT 297.750 266.215 301.300 266.715 ;
        RECT 0.000 264.980 6.000 266.030 ;
        RECT 295.300 265.165 301.300 266.215 ;
        RECT 0.000 264.280 3.555 264.980 ;
        RECT 297.750 264.265 301.300 265.165 ;
        RECT 0.000 259.970 3.555 260.670 ;
        RECT 297.750 260.155 301.300 260.655 ;
        RECT 0.000 258.920 6.000 259.970 ;
        RECT 295.300 259.105 301.300 260.155 ;
        RECT 0.000 258.220 3.555 258.920 ;
        RECT 297.750 258.205 301.300 259.105 ;
        RECT 0.000 253.910 3.555 254.610 ;
        RECT 297.750 254.095 301.300 254.595 ;
        RECT 0.000 252.860 6.000 253.910 ;
        RECT 295.300 253.045 301.300 254.095 ;
        RECT 0.000 252.160 3.555 252.860 ;
        RECT 297.750 252.145 301.300 253.045 ;
        RECT 0.000 247.850 3.555 248.550 ;
        RECT 297.750 248.035 301.300 248.535 ;
        RECT 0.000 246.800 6.000 247.850 ;
        RECT 295.300 246.985 301.300 248.035 ;
        RECT 0.000 246.100 3.555 246.800 ;
        RECT 297.750 246.085 301.300 246.985 ;
        RECT 0.000 241.790 3.555 242.490 ;
        RECT 297.750 241.975 301.300 242.475 ;
        RECT 0.000 240.740 6.000 241.790 ;
        RECT 295.300 240.925 301.300 241.975 ;
        RECT 0.000 240.040 3.555 240.740 ;
        RECT 297.750 240.025 301.300 240.925 ;
        RECT 0.000 235.730 3.555 236.430 ;
        RECT 297.750 235.915 301.300 236.415 ;
        RECT 0.000 234.680 6.000 235.730 ;
        RECT 295.300 234.865 301.300 235.915 ;
        RECT 0.000 233.980 3.555 234.680 ;
        RECT 297.750 233.965 301.300 234.865 ;
        RECT 0.000 229.670 3.555 230.370 ;
        RECT 297.750 229.855 301.300 230.355 ;
        RECT 0.000 228.620 6.000 229.670 ;
        RECT 295.300 228.805 301.300 229.855 ;
        RECT 0.000 227.920 3.555 228.620 ;
        RECT 297.750 227.905 301.300 228.805 ;
        RECT 0.000 223.610 3.555 224.310 ;
        RECT 297.750 223.795 301.300 224.295 ;
        RECT 0.000 222.560 6.000 223.610 ;
        RECT 295.300 222.745 301.300 223.795 ;
        RECT 0.000 221.860 3.555 222.560 ;
        RECT 297.750 221.845 301.300 222.745 ;
        RECT 0.000 217.550 3.555 218.250 ;
        RECT 297.750 217.735 301.300 218.235 ;
        RECT 0.000 216.500 6.000 217.550 ;
        RECT 295.300 216.685 301.300 217.735 ;
        RECT 0.000 215.800 3.555 216.500 ;
        RECT 297.750 215.785 301.300 216.685 ;
        RECT 0.000 211.490 3.555 212.190 ;
        RECT 297.750 211.675 301.300 212.175 ;
        RECT 0.000 210.440 6.000 211.490 ;
        RECT 295.300 210.625 301.300 211.675 ;
        RECT 0.000 209.740 3.555 210.440 ;
        RECT 297.750 209.725 301.300 210.625 ;
        RECT 0.000 205.430 3.555 206.130 ;
        RECT 297.750 205.615 301.300 206.115 ;
        RECT 0.000 204.380 6.000 205.430 ;
        RECT 295.300 204.565 301.300 205.615 ;
        RECT 0.000 203.680 3.555 204.380 ;
        RECT 297.750 203.665 301.300 204.565 ;
        RECT 0.000 199.370 3.555 200.070 ;
        RECT 297.750 199.555 301.300 200.055 ;
        RECT 0.000 198.320 6.000 199.370 ;
        RECT 295.300 198.505 301.300 199.555 ;
        RECT 0.000 197.620 3.555 198.320 ;
        RECT 297.750 197.605 301.300 198.505 ;
        RECT 0.000 193.310 3.555 194.010 ;
        RECT 297.750 193.495 301.300 193.995 ;
        RECT 0.000 192.260 6.000 193.310 ;
        RECT 295.300 192.445 301.300 193.495 ;
        RECT 0.000 191.560 3.555 192.260 ;
        RECT 297.750 191.545 301.300 192.445 ;
        RECT 0.000 187.250 3.555 187.950 ;
        RECT 297.750 187.435 301.300 187.935 ;
        RECT 0.000 186.200 6.000 187.250 ;
        RECT 295.300 186.385 301.300 187.435 ;
        RECT 0.000 185.500 3.555 186.200 ;
        RECT 297.750 185.485 301.300 186.385 ;
        RECT 0.000 181.190 3.555 181.890 ;
        RECT 297.750 181.375 301.300 181.875 ;
        RECT 0.000 180.140 6.000 181.190 ;
        RECT 295.300 180.325 301.300 181.375 ;
        RECT 0.000 179.440 3.555 180.140 ;
        RECT 297.750 179.425 301.300 180.325 ;
        RECT 0.000 175.130 3.555 175.830 ;
        RECT 297.750 175.315 301.300 175.815 ;
        RECT 0.000 174.080 6.000 175.130 ;
        RECT 295.300 174.265 301.300 175.315 ;
        RECT 0.000 173.380 3.555 174.080 ;
        RECT 297.750 173.365 301.300 174.265 ;
        RECT 0.000 169.070 3.555 169.770 ;
        RECT 297.750 169.255 301.300 169.755 ;
        RECT 0.000 168.020 6.000 169.070 ;
        RECT 295.300 168.205 301.300 169.255 ;
        RECT 0.000 167.320 3.555 168.020 ;
        RECT 297.750 167.305 301.300 168.205 ;
        RECT 0.000 163.010 3.555 163.710 ;
        RECT 297.750 163.195 301.300 163.695 ;
        RECT 0.000 161.960 6.000 163.010 ;
        RECT 295.300 162.145 301.300 163.195 ;
        RECT 0.000 161.260 3.555 161.960 ;
        RECT 297.750 161.245 301.300 162.145 ;
        RECT 0.000 156.950 3.555 157.650 ;
        RECT 297.750 157.135 301.300 157.635 ;
        RECT 0.000 155.900 6.000 156.950 ;
        RECT 295.300 156.085 301.300 157.135 ;
        RECT 0.000 155.200 3.555 155.900 ;
        RECT 297.750 155.185 301.300 156.085 ;
        RECT 0.000 150.890 3.555 151.590 ;
        RECT 297.750 151.075 301.300 151.575 ;
        RECT 0.000 149.840 6.000 150.890 ;
        RECT 295.300 150.025 301.300 151.075 ;
        RECT 0.000 149.140 3.555 149.840 ;
        RECT 297.750 149.125 301.300 150.025 ;
        RECT 0.000 144.830 3.555 145.530 ;
        RECT 297.750 145.015 301.300 145.515 ;
        RECT 0.000 143.780 6.000 144.830 ;
        RECT 295.300 143.965 301.300 145.015 ;
        RECT 0.000 143.080 3.555 143.780 ;
        RECT 297.750 143.065 301.300 143.965 ;
        RECT 0.000 138.770 3.555 139.470 ;
        RECT 297.750 138.955 301.300 139.455 ;
        RECT 0.000 137.720 6.000 138.770 ;
        RECT 295.300 137.905 301.300 138.955 ;
        RECT 0.000 137.020 3.555 137.720 ;
        RECT 297.750 137.005 301.300 137.905 ;
        RECT 0.000 132.710 3.555 133.410 ;
        RECT 297.750 132.895 301.300 133.395 ;
        RECT 0.000 131.660 6.000 132.710 ;
        RECT 295.300 131.845 301.300 132.895 ;
        RECT 0.000 130.960 3.555 131.660 ;
        RECT 297.750 130.945 301.300 131.845 ;
        RECT 0.000 126.650 3.555 127.350 ;
        RECT 297.755 127.190 301.300 127.335 ;
        RECT 297.750 126.835 301.300 127.190 ;
        RECT 0.000 125.600 6.000 126.650 ;
        RECT 295.300 125.785 301.300 126.835 ;
        RECT 0.000 124.900 3.555 125.600 ;
        RECT 297.750 124.885 301.300 125.785 ;
        RECT 0.000 120.590 3.555 121.290 ;
        RECT 297.755 121.080 301.300 121.275 ;
        RECT 297.750 120.775 301.300 121.080 ;
        RECT 0.000 119.540 6.000 120.590 ;
        RECT 295.300 119.725 301.300 120.775 ;
        RECT 0.000 118.840 3.555 119.540 ;
        RECT 297.750 118.825 301.300 119.725 ;
        RECT 0.010 114.115 6.000 114.360 ;
        RECT 0.000 113.660 6.000 114.115 ;
        RECT 295.300 113.660 301.300 114.360 ;
        RECT 0.000 113.025 3.555 113.660 ;
        RECT 297.750 113.025 301.300 113.660 ;
        RECT 0.000 111.350 6.000 113.025 ;
        RECT 0.010 111.345 6.000 111.350 ;
        RECT 295.300 111.345 301.300 113.025 ;
        RECT 0.000 93.825 3.545 93.830 ;
        RECT 297.750 93.825 301.300 93.830 ;
        RECT 0.000 86.895 6.000 93.825 ;
        RECT 0.010 86.890 6.000 86.895 ;
        RECT 295.300 86.890 301.300 93.825 ;
        RECT 295.300 86.830 295.500 86.890 ;
        RECT 0.000 72.855 0.700 72.860 ;
        RECT 297.755 72.855 301.300 72.860 ;
        RECT 0.000 71.265 6.000 72.855 ;
        RECT 295.300 71.265 301.300 72.855 ;
        RECT 0.000 69.355 3.555 71.265 ;
        RECT 297.755 70.860 301.300 71.265 ;
        RECT 297.750 69.355 301.300 70.860 ;
        RECT 0.000 47.950 6.000 57.210 ;
        RECT 295.300 47.950 301.300 57.210 ;
        RECT 297.750 38.225 301.300 38.230 ;
        RECT 0.000 33.615 6.000 38.225 ;
        RECT 295.300 33.615 301.300 38.225 ;
        RECT 0.000 23.645 6.000 25.465 ;
        RECT 295.300 23.645 301.300 25.465 ;
        RECT 0.000 23.315 3.565 23.645 ;
        RECT 297.745 23.315 301.300 23.645 ;
        RECT 0.000 21.325 3.555 23.315 ;
        RECT 297.750 21.325 301.300 23.315 ;
        RECT 0.000 19.810 6.000 21.325 ;
        RECT 295.300 19.810 301.300 21.325 ;
        RECT 0.000 13.195 0.700 13.200 ;
        RECT 0.000 11.965 6.000 13.195 ;
        RECT 295.300 11.965 301.300 13.195 ;
        RECT 0.000 9.985 3.545 11.965 ;
        RECT 297.805 9.985 301.300 11.965 ;
        RECT 0.000 8.740 6.000 9.985 ;
        RECT 295.300 8.750 301.300 9.985 ;
        RECT 295.300 8.745 298.065 8.750 ;
        RECT 16.245 0.000 19.745 3.260 ;
        RECT 33.045 0.000 36.545 3.260 ;
        RECT 54.045 0.000 57.545 3.260 ;
        RECT 70.845 0.000 74.345 3.260 ;
        RECT 109.630 0.000 113.130 3.260 ;
        RECT 115.575 0.000 119.075 3.260 ;
        RECT 121.905 0.000 125.405 3.260 ;
        RECT 133.095 0.000 136.595 3.260 ;
        RECT 144.315 0.000 147.815 3.260 ;
        RECT 152.715 0.000 156.215 3.260 ;
        RECT 161.115 0.000 164.615 3.260 ;
        RECT 179.315 0.000 182.815 3.260 ;
        RECT 183.670 0.000 187.170 3.260 ;
        RECT 223.760 0.000 227.260 3.260 ;
        RECT 240.560 0.000 244.060 3.260 ;
        RECT 261.560 0.000 265.060 3.260 ;
        RECT 278.360 0.000 281.860 3.260 ;
    END
  END VSS
  PIN WEN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 288.510 5.985 289.140 5.990 ;
        RECT 288.510 5.955 289.420 5.985 ;
        RECT 288.510 5.695 290.025 5.955 ;
        RECT 288.510 5.685 289.420 5.695 ;
        RECT 288.510 5.650 289.140 5.685 ;
      LAYER Metal2 ;
        RECT 288.430 0.000 289.215 5.995 ;
    END
  END WEN[7]
  PIN WEN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 253.790 5.985 254.350 5.995 ;
        RECT 253.285 5.965 254.350 5.985 ;
        RECT 253.185 5.705 254.355 5.965 ;
        RECT 253.285 5.695 254.350 5.705 ;
        RECT 253.285 5.645 253.915 5.695 ;
      LAYER Metal2 ;
        RECT 253.205 0.000 253.985 6.000 ;
    END
  END WEN[6]
  PIN WEN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 249.780 5.950 250.340 5.980 ;
        RECT 250.710 5.950 251.340 5.985 ;
        RECT 249.775 5.690 251.340 5.950 ;
        RECT 249.780 5.680 250.340 5.690 ;
        RECT 250.710 5.645 251.340 5.690 ;
      LAYER Metal2 ;
        RECT 250.630 0.000 251.410 6.000 ;
    END
  END WEN[5]
  PIN WEN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 214.710 5.960 215.270 5.990 ;
        RECT 214.105 5.950 215.275 5.960 ;
        RECT 214.105 5.940 216.880 5.950 ;
        RECT 214.105 5.700 217.110 5.940 ;
        RECT 214.320 5.690 217.110 5.700 ;
        RECT 216.480 5.600 217.110 5.690 ;
        RECT 216.525 5.505 216.880 5.600 ;
      LAYER Metal2 ;
        RECT 216.400 0.000 217.185 5.955 ;
    END
  END WEN[4]
  PIN WEN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 81.990 5.975 82.620 5.990 ;
        RECT 83.305 5.975 83.865 5.980 ;
        RECT 81.950 5.950 84.110 5.975 ;
        RECT 81.950 5.690 84.470 5.950 ;
        RECT 81.950 5.670 84.110 5.690 ;
        RECT 81.990 5.650 82.620 5.670 ;
      LAYER Metal2 ;
        RECT 81.910 0.000 82.695 6.000 ;
    END
  END WEN[3]
  PIN WEN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 45.915 5.940 46.545 5.990 ;
        RECT 48.235 5.960 48.795 5.990 ;
        RECT 47.630 5.940 48.800 5.960 ;
        RECT 45.915 5.700 48.800 5.940 ;
        RECT 45.915 5.690 48.795 5.700 ;
        RECT 45.915 5.665 48.390 5.690 ;
        RECT 45.915 5.650 46.545 5.665 ;
      LAYER Metal2 ;
        RECT 45.685 5.650 46.545 5.990 ;
        RECT 45.685 0.000 46.470 5.650 ;
    END
  END WEN[2]
  PIN WEN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 44.190 5.980 44.820 5.990 ;
        RECT 44.190 5.950 45.035 5.980 ;
        RECT 44.190 5.690 45.640 5.950 ;
        RECT 44.190 5.680 45.035 5.690 ;
        RECT 44.190 5.665 44.945 5.680 ;
        RECT 44.190 5.650 44.820 5.665 ;
      LAYER Metal2 ;
        RECT 44.110 0.000 44.895 5.995 ;
    END
  END WEN[1]
  PIN WEN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.800 5.650 10.850 6.000 ;
        RECT 10.215 5.645 10.845 5.650 ;
      LAYER Metal2 ;
        RECT 10.215 5.980 10.845 5.985 ;
        RECT 10.085 0.000 10.870 5.980 ;
    END
  END WEN[0]
  OBS
      LAYER Nwell ;
        RECT 6.305 6.000 295.010 315.890 ;
      LAYER Metal1 ;
        RECT 6.000 6.000 295.300 315.890 ;
      LAYER Metal2 ;
        RECT 6.000 6.000 295.300 315.890 ;
      LAYER Metal3 ;
        RECT 6.000 86.350 295.300 315.890 ;
        RECT 6.000 85.600 295.500 86.350 ;
        RECT 6.000 85.125 295.300 85.600 ;
        RECT 6.000 84.370 295.500 85.125 ;
        RECT 6.000 83.900 295.300 84.370 ;
        RECT 6.000 83.145 295.500 83.900 ;
        RECT 6.000 82.675 295.300 83.145 ;
        RECT 6.000 81.920 295.500 82.675 ;
        RECT 6.000 6.000 295.300 81.920 ;
  END
END gf180mcu_ocd_ip_sram__sram512x8m8wm1
END LIBRARY

