magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< polysilicon >>
rect -14 943 41 975
rect -14 -33 41 0
use nmos_5p04310591302099_512x8m81  nmos_5p04310591302099_512x8m81_0
timestamp 1763476864
transform 1 0 -14 0 1 0
box -88 -44 144 987
<< end >>
