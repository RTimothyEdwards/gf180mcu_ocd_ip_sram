magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal1 >>
rect -113 1146 113 1155
rect -113 -1146 -105 1146
rect 105 -1146 113 1146
rect -113 -1155 113 -1146
<< via1 >>
rect -105 -1146 105 1146
<< metal2 >>
rect -113 1146 113 1155
rect -113 -1146 -105 1146
rect 105 -1146 113 1146
rect -113 -1155 113 -1146
<< end >>
