magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< error_s >>
rect 19225 45914 19230 45919
rect 19271 25190 19276 45914
rect 39909 25190 39915 45919
rect 19209 24246 19236 24302
rect 19225 24240 19230 24246
rect 19265 23908 19292 24246
<< psubdiff >>
rect 18967 25183 20040 46016
rect 39151 25183 40172 46326
rect 59602 2309 59871 46323
<< metal1 >>
rect 0 2187 700 46294
<< metal2 >>
rect 296 2187 996 46301
<< metal3 >>
rect 296 2722 997 2791
rect 296 1905 996 2722
use M1_PSUB4310591302043_3v256x8m81  M1_PSUB4310591302043_3v256x8m81_0
timestamp 1763766357
transform -1 0 59970 0 1 46009
box 171 -29 59921 289
use M1_PSUB4310591302043_3v256x8m81  M1_PSUB4310591302043_3v256x8m81_1
timestamp 1763766357
transform -1 0 59970 0 1 2339
box 171 -29 59921 289
use M1_PSUB4310591302044_3v256x8m81  M1_PSUB4310591302044_3v256x8m81_0
timestamp 1763766357
transform 1 0 59631 0 1 798
box -29 1830 240 45182
use M1_PSUB4310591302044_3v256x8m81  M1_PSUB4310591302044_3v256x8m81_1
timestamp 1763766357
transform 1 0 18997 0 1 798
box -29 1830 240 45182
use M1_PSUB4310591302044_3v256x8m81  M1_PSUB4310591302044_3v256x8m81_2
timestamp 1763766357
transform 1 0 39932 0 1 798
box -29 1830 240 45182
use M1_PSUB4310591302044_3v256x8m81  M1_PSUB4310591302044_3v256x8m81_3
timestamp 1763766357
transform 1 0 78 0 1 798
box -29 1830 240 45182
use M1_PSUB4310591302045_3v256x8m81  M1_PSUB4310591302045_3v256x8m81_0
timestamp 1763766357
transform 1 0 39286 0 1 25213
box -29 -29 589 20707
use M1_PSUB4310591302045_3v256x8m81  M1_PSUB4310591302045_3v256x8m81_1
timestamp 1763766357
transform 1 0 19294 0 1 25213
box -29 -29 589 20707
use M1_PSUB4310591302046_3v256x8m81  M1_PSUB4310591302046_3v256x8m81_0
timestamp 1763766357
transform 1 0 19294 0 1 23937
box -29 -29 20539 309
<< labels >>
flabel metal3 s 646 2029 646 2029 0 FreeSans 313 0 0 0 VDD
port 1 nsew
<< properties >>
string path 4.620 11.160 4.620 0.000 
<< end >>
