magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal2 >>
rect -35 628 35 635
rect -35 -628 -28 628
rect 28 -628 35 628
rect -35 -635 35 -628
<< via2 >>
rect -28 -628 28 628
<< metal3 >>
rect -35 628 35 635
rect -35 -628 -28 628
rect 28 -628 35 628
rect -35 -635 35 -628
<< end >>
