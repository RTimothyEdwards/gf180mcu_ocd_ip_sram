magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< metal1 >>
rect -413 26 413 46
rect -413 -26 -395 26
rect 395 -26 413 26
rect -413 -46 413 -26
<< via1 >>
rect -395 -26 395 26
<< metal2 >>
rect -414 26 414 46
rect -414 -26 -395 26
rect 395 -26 414 26
rect -414 -46 414 -26
<< end >>
