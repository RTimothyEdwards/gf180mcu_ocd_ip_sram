magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< nwell >>
rect 798 5267 1239 5500
rect -134 3584 -130 5026
rect 217 4720 1239 5267
rect 265 4380 1239 4720
rect 798 3571 1239 4380
rect 1332 1103 1824 1115
rect 208 959 1824 1103
rect -156 406 1824 959
rect 207 405 806 406
rect 1383 405 1824 406
rect 208 348 806 405
rect 1384 -35 1824 405
<< nmos >>
rect 522 5417 578 5524
<< pmos >>
rect 451 5030 507 5169
rect 614 5030 670 5169
<< ndiff >>
rect 406 5476 522 5524
rect 406 5430 437 5476
rect 483 5430 522 5476
rect 406 5417 522 5430
rect 578 5476 684 5524
rect 578 5430 621 5476
rect 667 5430 684 5476
rect 578 5417 684 5430
<< pdiff >>
rect 340 5095 451 5169
rect 340 5049 357 5095
rect 403 5049 451 5095
rect 340 5030 451 5049
rect 507 5095 614 5169
rect 507 5049 539 5095
rect 585 5049 614 5095
rect 507 5030 614 5049
rect 670 5095 781 5169
rect 670 5049 719 5095
rect 765 5049 781 5095
rect 670 5030 781 5049
<< ndiffc >>
rect 437 5430 483 5476
rect 621 5430 667 5476
<< pdiffc >>
rect 357 5049 403 5095
rect 539 5049 585 5095
rect 719 5049 765 5095
<< polysilicon >>
rect 522 5524 578 5575
rect 522 5316 578 5417
rect 451 5218 670 5316
rect 451 5169 507 5218
rect 614 5169 670 5218
rect 451 4980 507 5030
rect 614 4980 670 5030
rect 497 4708 633 4855
rect 357 4666 727 4708
rect 357 4344 413 4666
rect 671 4344 727 4666
rect 44 2755 100 3640
rect 997 3564 1053 3635
rect 908 3469 1053 3564
rect 997 2878 1053 3469
rect 357 1671 727 1735
rect 966 1514 1050 1581
rect 976 1510 1032 1514
rect 44 1405 100 1424
rect 976 1276 1032 1342
rect 976 1234 1193 1276
rect 471 1084 527 1223
rect 976 1178 1032 1234
rect 1136 1176 1192 1234
rect 401 1041 617 1084
rect 401 771 457 858
rect 767 786 1197 828
rect 387 730 471 771
rect 387 688 1037 730
rect 981 632 1037 688
rect 1141 635 1197 786
rect 1533 738 1589 1280
rect 419 370 475 425
rect 194 328 475 370
rect 194 327 329 328
rect 419 273 475 328
rect 579 272 635 430
rect 981 407 1036 478
rect 981 364 1179 407
rect 795 267 1019 309
rect 963 234 1019 267
rect 1123 230 1179 364
<< metal1 >>
rect 248 6117 1446 6185
rect 248 5971 1446 6038
rect 31 5796 1446 5892
rect 114 5647 1106 5714
rect 413 5536 825 5587
rect 413 5476 494 5536
rect -32 4761 16 5469
rect 413 5430 437 5476
rect 483 5430 494 5476
rect 413 5424 494 5430
rect 562 5476 678 5488
rect 562 5430 621 5476
rect 667 5430 678 5476
rect 562 5387 678 5430
rect 326 5222 507 5315
rect 562 5163 612 5387
rect 346 5095 414 5154
rect 346 5049 357 5095
rect 403 5049 414 5095
rect 346 5036 414 5049
rect 531 5095 612 5163
rect 531 5049 539 5095
rect 585 5049 612 5095
rect 531 5036 612 5049
rect 363 4725 414 5036
rect 562 4781 612 5036
rect 694 5095 775 5163
rect 694 5082 719 5095
rect 694 5049 718 5082
rect 765 5049 775 5095
rect 694 5036 775 5049
rect 694 4725 744 5036
rect 1081 4727 1128 5445
rect 363 4673 744 4725
rect 278 4276 335 4404
rect 588 4274 645 4402
rect 116 3558 197 3863
rect 429 3558 511 3863
rect 923 3760 973 3863
rect 743 3676 973 3760
rect 116 3474 877 3558
rect -31 2677 19 3333
rect 116 2688 197 3474
rect 274 2797 334 3319
rect 429 2765 511 3474
rect 923 3358 973 3676
rect 1396 3366 1508 5422
rect 591 2816 651 3329
rect 754 3274 973 3358
rect 754 2786 814 3274
rect 923 2775 973 3274
rect 1057 1817 1508 3366
rect 432 1659 634 1726
rect 251 1519 1512 1603
rect 251 1389 332 1519
rect 37 1305 332 1389
rect 577 1125 627 1342
rect 486 1073 836 1125
rect 486 904 536 1073
rect 158 689 443 765
rect 135 307 286 391
rect 340 375 391 500
rect 340 323 590 375
rect 0 62 46 198
rect 340 172 391 323
rect 490 62 540 170
rect 0 10 540 62
rect 684 62 734 536
rect 785 273 836 1073
rect 889 828 970 1098
rect 900 827 966 828
rect 1045 772 1127 1433
rect 1202 828 1283 998
rect 1045 688 1283 772
rect 888 62 934 571
rect 684 10 934 62
rect 1081 13 1128 556
rect 1202 101 1283 688
rect 1458 624 1512 1519
rect 1648 1294 1725 1510
rect 1618 649 1707 865
rect 1081 -38 1590 13
<< metal2 >>
rect 277 3133 343 6185
rect 558 6044 621 6304
rect 558 5961 658 6044
rect 436 1663 501 5892
rect 592 3133 658 5961
rect 803 5579 869 6415
rect 1052 6117 1115 6264
rect 1463 5971 1525 6301
rect 752 5511 869 5579
rect 752 5355 818 5511
rect 767 221 833 1349
rect 485 153 833 221
<< metal3 >>
rect -32 3630 1719 5535
rect -32 1048 1719 3430
rect -32 441 1719 943
use M1_NWELL08_512x8m81  M1_NWELL08_512x8m81_0
timestamp 1763476864
transform 1 0 0 0 1 742
box -154 -216 154 216
use M1_NWELL4310591302032_512x8m81  M1_NWELL4310591302032_512x8m81_0
timestamp 1763476864
transform 1 0 1021 0 1 5408
box -126 -85 127 87
use M1_PACTIVE4310591302027_512x8m81  M1_PACTIVE4310591302027_512x8m81_0
timestamp 1763476864
transform 1 0 23 0 1 174
box -36 -62 36 62
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1763476864
transform 1 0 473 0 1 1699
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1763476864
transform 1 0 810 0 1 296
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_2
timestamp 1763476864
transform 1 0 1559 0 1 -14
box -36 -36 36 36
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_3
timestamp 1763476864
transform 1 0 1008 0 1 1551
box -36 -36 36 36
use M1_PSUB$$45111340_512x8m81  M1_PSUB$$45111340_512x8m81_0
timestamp 1763476864
transform 1 0 0 0 1 1183
box -56 -58 56 58
use M1_PSUB$$46892076_512x8m81  M1_PSUB$$46892076_512x8m81_0
timestamp 1763476864
transform 1 0 1446 0 1 3657
box -56 -1771 56 1771
use M1_PSUB$$46893100_512x8m81  M1_PSUB$$46893100_512x8m81_0
timestamp 1763476864
transform 1 0 1335 0 1 2629
box -56 -742 56 743
use M2_M1$$43375660_R90_512x8m81  M2_M1$$43375660_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 73 1 0 1180
box -46 -119 46 119
use M2_M1$$46894124_512x8m81  M2_M1$$46894124_512x8m81_0
timestamp 1763476864
transform 1 0 469 0 1 5846
box -44 -46 45 46
use M3_M2$$43368492_R90_512x8m81  M3_M2$$43368492_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 73 1 0 1180
box -46 -119 46 119
use M3_M2$$46895148_512x8m81  M3_M2$$46895148_512x8m81_0
timestamp 1763476864
transform 1 0 469 0 1 5846
box -45 -46 45 46
use nmos_1p2$$46563372_512x8m81  nmos_1p2$$46563372_512x8m81_0
timestamp 1763476864
transform 1 0 990 0 -1 1469
box -102 -44 130 133
use nmos_1p2$$46563372_512x8m81  nmos_1p2$$46563372_512x8m81_1
timestamp 1763476864
transform 1 0 485 0 1 1264
box -102 -44 130 133
use nmos_1p2$$46883884_512x8m81  nmos_1p2$$46883884_512x8m81_0
timestamp 1763476864
transform 1 0 685 0 1 1777
box -102 -44 130 1102
use nmos_1p2$$46883884_512x8m81  nmos_1p2$$46883884_512x8m81_1
timestamp 1763476864
transform 1 0 1011 0 1 1777
box -102 -44 130 1102
use nmos_1p2$$46883884_512x8m81  nmos_1p2$$46883884_512x8m81_2
timestamp 1763476864
transform 1 0 371 0 1 1777
box -102 -44 130 1102
use nmos_1p2$$46884908_512x8m81  nmos_1p2$$46884908_512x8m81_0
timestamp 1763476864
transform 1 0 58 0 1 1460
box -102 -44 130 1314
use nmos_5p04310591302010_512x8m81  nmos_5p04310591302010_512x8m81_0
timestamp 1763476864
transform 1 0 1533 0 -1 1529
box -88 -44 144 255
use nmos_5p04310591302011_512x8m81  nmos_5p04310591302011_512x8m81_0
timestamp 1763476864
transform 1 0 447 0 -1 250
box -116 -44 276 133
use nmos_5p04310591302011_512x8m81  nmos_5p04310591302011_512x8m81_1
timestamp 1763476864
transform 1 0 991 0 1 101
box -116 -44 276 133
use pmos_1p2$$46273580_512x8m81  pmos_1p2$$46273580_512x8m81_0
timestamp 1763476864
transform 1 0 443 0 -1 1004
box -216 -86 348 192
use pmos_1p2$$46273580_512x8m81  pmos_1p2$$46273580_512x8m81_1
timestamp 1763476864
transform 1 0 1018 0 -1 1139
box -216 -86 348 192
use pmos_1p2$$46885932_512x8m81  pmos_1p2$$46885932_512x8m81_0
timestamp 1763476864
transform 1 0 1023 0 1 504
box -216 -86 348 175
use pmos_1p2$$46887980_512x8m81  pmos_1p2$$46887980_512x8m81_0
timestamp 1763476864
transform 1 0 58 0 1 3670
box -188 -86 216 1356
use pmos_1p2$$46889004_512x8m81  pmos_1p2$$46889004_512x8m81_0
timestamp 1763476864
transform 1 0 371 0 1 3670
box -188 -86 216 721
use pmos_1p2$$46889004_512x8m81  pmos_1p2$$46889004_512x8m81_1
timestamp 1763476864
transform 1 0 685 0 1 3670
box -188 -86 216 721
use pmos_5p0431059130201_512x8m81  pmos_5p0431059130201_512x8m81_0
timestamp 1763476864
transform 1 0 1533 0 1 63
box -174 -86 230 721
use pmos_5p0431059130206_512x8m81  pmos_5p0431059130206_512x8m81_0
timestamp 1763476864
transform 1 0 447 0 1 447
box -202 -86 362 175
use pmos_5p0431059130209_512x8m81  pmos_5p0431059130209_512x8m81_0
timestamp 1763476864
transform 1 0 997 0 1 3670
box -174 -86 230 1144
use po_m1_512x8m81  po_m1_512x8m81_0
timestamp 1763476864
transform -1 0 638 0 -1 396
box -21 0 113 95
use po_m1_512x8m81  po_m1_512x8m81_1
timestamp 1763476864
transform 1 0 519 0 -1 4854
box -21 0 113 95
use po_m1_512x8m81  po_m1_512x8m81_2
timestamp 1763476864
transform 1 0 356 0 1 688
box -21 0 113 95
use po_m1_512x8m81  po_m1_512x8m81_3
timestamp 1763476864
transform 1 0 32 0 1 1313
box -21 0 113 95
use po_m1_R90_512x8m81  po_m1_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 897 1 0 3469
box 0 -21 95 113
use po_m1_R90_512x8m81  po_m1_R90_512x8m81_1
timestamp 1763476864
transform 0 -1 847 1 0 786
box 0 -21 95 113
use po_m1_R270_512x8m81  po_m1_R270_512x8m81_0
timestamp 1763476864
transform 0 1 214 -1 0 396
box 0 -21 95 114
use po_m1_R270_512x8m81  po_m1_R270_512x8m81_1
timestamp 1763476864
transform 0 1 436 -1 0 5320
box 0 -21 95 114
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_0
timestamp 1763476864
transform -1 0 565 0 -1 676
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_1
timestamp 1763476864
transform -1 0 702 0 -1 920
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_2
timestamp 1763476864
transform -1 0 965 0 -1 920
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_3
timestamp 1763476864
transform 1 0 -32 0 1 2466
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_4
timestamp 1763476864
transform 1 0 1057 0 1 1824
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_5
timestamp 1763476864
transform 1 0 -22 0 1 3129
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_6
timestamp 1763476864
transform 1 0 1057 0 1 3129
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_7
timestamp 1763476864
transform 1 0 1057 0 1 2466
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_8
timestamp 1763476864
transform 1 0 -32 0 1 628
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_9
timestamp 1763476864
transform 1 0 402 0 1 1228
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_10
timestamp 1763476864
transform 1 0 1714 0 1 650
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_11
timestamp 1763476864
transform 1 0 1066 0 1 3826
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_12
timestamp 1763476864
transform 1 0 -32 0 1 3826
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_13
timestamp 1763476864
transform 1 0 1066 0 1 4869
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_14
timestamp 1763476864
transform 1 0 -32 0 1 5265
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_15
timestamp 1763476864
transform 1 0 -32 0 1 4846
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_16
timestamp 1763476864
transform 1 0 1714 0 1 1295
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_17
timestamp 1763476864
transform 1 0 905 0 1 1228
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_18
timestamp 1763476864
transform 1 0 -32 0 1 1824
box -9 0 73 215
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_19
timestamp 1763476864
transform 1 0 723 0 1 4939
box -9 0 73 215
use via1_2_x2_R90_512x8m81  via1_2_x2_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 390 1 0 854
box -9 0 73 215
use via1_2_x2_R90_512x8m81  via1_2_x2_R90_512x8m81_1
timestamp 1763476864
transform 0 -1 1128 1 0 5376
box -9 0 73 215
use via1_512x8m81  via1_512x8m81_0
timestamp 1763476864
transform 1 0 485 0 1 139
box 0 0 65 92
use via1_512x8m81  via1_512x8m81_1
timestamp 1763476864
transform 1 0 436 0 1 5222
box 0 0 65 92
use via1_R90_512x8m81  via1_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 522 1 0 1659
box 0 0 65 89
use via1_x2_512x8m81  via1_x2_512x8m81_0
timestamp 1763476864
transform -1 0 1268 0 -1 1050
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_1
timestamp 1763476864
transform 1 0 595 0 1 4387
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_2
timestamp 1763476864
transform 1 0 277 0 1 4387
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_3
timestamp 1763476864
transform 1 0 753 0 1 5355
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_4
timestamp 1763476864
transform 1 0 280 0 1 3133
box -8 0 72 222
use via1_x2_512x8m81  via1_x2_512x8m81_5
timestamp 1763476864
transform 1 0 595 0 1 3133
box -8 0 72 222
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_0
timestamp 1763476864
transform 0 -1 1610 1 0 5971
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_1
timestamp 1763476864
transform 0 -1 1190 1 0 6117
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_2
timestamp 1763476864
transform 0 -1 744 1 0 5971
box -8 0 72 215
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_3
timestamp 1763476864
transform 0 -1 448 1 0 6117
box -8 0 72 215
use via2_x2_512x8m81  via2_x2_512x8m81_0
timestamp 1763476864
transform -1 0 1268 0 -1 920
box -9 0 74 222
use via2_x2_512x8m81  via2_x2_512x8m81_1
timestamp 1763476864
transform 1 0 768 0 1 1127
box -9 0 74 222
<< labels >>
rlabel metal3 s 1089 2256 1089 2256 4 vss
port 1 nsew
rlabel metal3 s 1040 4168 1040 4168 4 vdd
port 2 nsew
rlabel metal3 s 935 642 935 642 4 vdd
port 2 nsew
rlabel metal2 s 304 5597 304 5597 4 d
port 3 nsew
rlabel metal1 s 263 355 263 355 4 datain
port 5 nsew
rlabel metal1 s 735 5854 735 5854 4 wep
port 6 nsew
rlabel metal1 s 399 739 399 739 4 men
port 7 nsew
rlabel metal1 s 877 6158 877 6158 4 d
port 3 nsew
rlabel metal1 s 975 6015 975 6015 4 db
port 4 nsew
rlabel metal2 s 829 5737 829 5737 4 vss
port 1 nsew
rlabel metal2 s 618 5597 618 5597 4 db
port 4 nsew
<< end >>
