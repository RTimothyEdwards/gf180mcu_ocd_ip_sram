magic
tech gf180mcuD
magscale 1 10
timestamp 1765899468
<< nwell >>
rect 20780 43711 38804 43962
rect 20780 43679 27872 43711
rect 20780 43472 22995 43679
rect 24681 43473 27872 43679
rect 24682 43472 27872 43473
rect 31637 43661 38804 43711
rect 31637 43472 34834 43661
rect 36598 43472 38804 43661
<< psubdiff >>
rect 19420 22003 40130 22342
<< metal1 >>
rect 197 44088 60063 44788
rect 197 897 897 44088
rect 18028 43115 18537 44088
rect 19324 23589 20437 44088
rect 23958 43372 24509 44088
rect 28043 43372 28413 44088
rect 30616 43372 31194 44088
rect 35068 43242 35639 44088
rect 19170 23284 20437 23589
rect 38969 23284 40415 44088
rect 40953 43115 41462 44088
rect 19170 22336 19479 23284
rect 40106 22336 40415 23284
rect 59363 22993 60063 44088
rect 58864 22871 60063 22993
rect 19170 22009 40415 22336
rect 1760 1130 2170 1200
rect 18740 1198 19049 21558
rect 19170 1302 19479 22009
rect 34809 4205 35009 4237
rect 34974 3400 36262 3448
rect 40106 1302 40415 22009
rect 8934 1133 8989 1174
rect 9198 1133 9678 1188
rect 16390 1134 16822 1195
rect 19170 897 40415 1302
rect 40536 1255 40845 21558
rect 58183 20528 58798 20580
rect 42824 1138 43436 1190
rect 59363 897 60063 22871
rect 197 896 40501 897
rect 40936 896 60063 897
rect 197 197 60063 896
<< metal2 >>
rect 197 44560 60063 44788
rect 494 43726 59766 44426
rect 494 3963 1194 43726
rect 18029 17339 18537 43532
rect 18627 17422 18937 43726
rect 19170 43475 19479 43478
rect 19170 43322 20812 43475
rect 19170 42249 19479 43322
rect 20964 43242 21374 43726
rect 21538 43242 23021 43726
rect 24589 43242 25490 43726
rect 27267 43372 27732 43726
rect 34152 43242 34993 43726
rect 36558 43242 38047 43726
rect 38209 43242 38619 43726
rect 38759 43334 40161 43479
rect 19170 42110 20849 42249
rect 38759 42122 40161 42237
rect 19170 41037 19479 42110
rect 19170 40898 20849 41037
rect 38759 40910 40161 41025
rect 19170 39825 19479 40898
rect 19170 39686 20849 39825
rect 38759 39698 40161 39813
rect 19170 38613 19479 39686
rect 19170 38474 20849 38613
rect 38759 38486 40161 38601
rect 19170 37401 19479 38474
rect 19170 37262 20849 37401
rect 38759 37274 40161 37389
rect 19170 36189 19479 37262
rect 19170 36050 20849 36189
rect 38759 36062 40161 36177
rect 19170 34977 19479 36050
rect 19170 34838 20849 34977
rect 38759 34850 40161 34965
rect 19170 33765 19479 34838
rect 19170 33626 20849 33765
rect 38759 33638 40161 33753
rect 19170 32553 19479 33626
rect 19170 32414 20849 32553
rect 38759 32426 40161 32541
rect 19170 31341 19479 32414
rect 19170 31202 20849 31341
rect 38759 31214 40161 31329
rect 19170 30129 19479 31202
rect 19170 29990 20849 30129
rect 38759 30002 40161 30117
rect 19170 28917 19479 29990
rect 19170 28778 20849 28917
rect 38759 28790 40161 28905
rect 19170 27705 19479 28778
rect 19170 27566 20849 27705
rect 38759 27578 40161 27693
rect 19170 26493 19479 27566
rect 19170 26354 20849 26493
rect 38759 26366 40161 26481
rect 19170 25281 19479 26354
rect 19170 25142 20849 25281
rect 38759 25154 40161 25269
rect 19170 24069 19479 25142
rect 19170 23930 20849 24069
rect 38759 23942 40161 24057
rect 19170 20772 19479 23930
rect 25804 23145 26420 23750
rect 29030 23127 29185 23362
rect 29295 23230 29450 23362
rect 27017 22967 29185 23127
rect 27017 22956 27171 22967
rect 22150 22795 27171 22956
rect 29295 22892 29450 23040
rect 22150 21439 22305 22795
rect 27353 22732 29450 22892
rect 27353 22714 27508 22732
rect 22399 22555 27508 22714
rect 29559 22658 29714 23362
rect 22399 21423 22554 22555
rect 27828 22497 29714 22658
rect 27828 22487 27983 22497
rect 26810 22327 27983 22487
rect 29822 22422 29977 23354
rect 26810 22238 26966 22327
rect 26040 22079 26966 22238
rect 28074 22263 29977 22422
rect 28074 22233 28229 22263
rect 26040 21447 26196 22079
rect 27049 22073 28229 22233
rect 30088 22188 30243 23362
rect 27049 22004 27204 22073
rect 26289 21843 27204 22004
rect 28320 22028 30243 22188
rect 28320 21998 28475 22028
rect 26289 21439 26444 21843
rect 27315 21838 28475 21998
rect 30351 21953 30506 23354
rect 31859 23184 32014 23362
rect 27315 21447 27470 21838
rect 28566 21793 30506 21953
rect 31252 23024 32014 23184
rect 28566 21752 28721 21793
rect 27562 21592 28721 21752
rect 31252 21598 31406 23024
rect 32123 22949 32278 23362
rect 31497 22789 32278 22949
rect 32387 23071 32543 23362
rect 32387 22912 32550 23071
rect 31497 21598 31653 22789
rect 32395 21598 32550 22912
rect 32652 22837 32807 23354
rect 32641 22676 32807 22837
rect 27562 21522 27717 21592
rect 32641 21589 32796 22676
rect 32918 22480 33073 23354
rect 33181 22714 33336 23362
rect 33445 22949 33600 23362
rect 33709 23184 33865 23362
rect 33709 23024 35084 23184
rect 33445 22789 34838 22949
rect 33181 22555 33940 22714
rect 32918 22319 33694 22480
rect 33539 21589 33694 22319
rect 33785 21598 33940 22555
rect 34682 21598 34838 22789
rect 34928 21598 35084 23024
rect 18803 17262 18897 17422
rect 17289 11780 17389 15565
rect 17480 12018 17580 15808
rect 17650 12257 17750 16050
rect 17826 12494 17926 16289
rect 18004 12732 18104 16523
rect 18178 12970 18278 16757
rect 18353 13208 18453 17010
rect 18544 13446 18644 17233
rect 740 3928 1194 3963
rect 494 2844 1194 3928
rect 1766 3293 1831 3524
rect 739 2757 1194 2844
rect 494 197 1194 2757
rect 1304 3216 1831 3293
rect 2389 3402 2455 3517
rect 8443 3404 8509 3548
rect 2389 3359 2459 3402
rect 2389 3276 2517 3359
rect 2394 3275 2517 3276
rect 1304 3215 1797 3216
rect 1304 0 1461 3215
rect 2017 0 2174 1196
rect 2451 1156 2517 3275
rect 8309 3338 8509 3404
rect 2451 1090 2883 1156
rect 2817 849 2883 1090
rect 8309 945 8375 3338
rect 9055 3326 9120 3554
rect 8835 3261 9120 3326
rect 9537 3337 9602 3581
rect 10155 3428 10221 3579
rect 10155 3362 10316 3428
rect 9537 3280 9803 3337
rect 8835 1321 8900 3261
rect 8643 1256 8900 1321
rect 8643 1058 8708 1256
rect 8168 879 8375 945
rect 2766 0 2922 849
rect 8168 840 8234 879
rect 8073 711 8234 840
rect 8636 834 8708 1058
rect 8073 0 8229 711
rect 8544 0 8701 834
rect 8822 0 8979 1199
rect 9137 0 9294 1198
rect 9746 1085 9803 3280
rect 10250 1090 10316 3362
rect 16209 3287 16275 3545
rect 15595 3221 16275 3287
rect 16818 3293 16883 3523
rect 17139 3293 17200 3294
rect 9519 1028 9803 1085
rect 9519 832 9576 1028
rect 9992 1024 10316 1090
rect 9992 832 10058 1024
rect 9417 744 9576 832
rect 9417 0 9574 744
rect 9888 742 10058 832
rect 15596 826 15663 3221
rect 16818 3215 17200 3293
rect 9888 0 10045 742
rect 15595 0 15752 826
rect 16382 0 16539 1200
rect 17139 970 17200 3215
rect 19170 1762 19479 20672
rect 34970 4210 35028 6046
rect 36225 3395 36283 6711
rect 16656 909 17200 970
rect 16656 0 16813 909
rect 19555 0 19712 2126
rect 20304 1525 20394 2151
rect 20472 1861 20563 2151
rect 20472 1696 20950 1861
rect 20304 290 20461 1525
rect 20793 0 20950 1696
rect 21601 0 21758 2455
rect 22786 0 22943 2455
rect 23970 0 24126 2455
rect 28411 0 28568 2088
rect 35239 0 35396 3189
rect 37640 2011 38968 2168
rect 37640 0 37797 2011
rect 39046 1855 39137 2131
rect 38091 1699 39137 1855
rect 38091 0 38248 1699
rect 39216 1517 39306 2131
rect 38614 1360 39306 1517
rect 38614 0 38771 1360
rect 39385 0 39542 2349
rect 40106 1766 40415 21558
rect 40536 1766 40845 43726
rect 40953 17390 41461 43598
rect 59089 43062 59766 43726
rect 59088 22087 59766 43062
rect 59066 7916 59766 22087
rect 59066 7458 59767 7916
rect 42832 3293 42897 3526
rect 42451 3215 42897 3293
rect 43450 3359 43516 3515
rect 49509 3405 49566 3526
rect 43450 3275 43638 3359
rect 42451 871 42525 3215
rect 43280 1180 43437 1191
rect 43280 1128 43305 1180
rect 43413 1128 43437 1180
rect 42451 870 42788 871
rect 42451 797 42969 870
rect 42812 0 42969 797
rect 43280 0 43437 1128
rect 43572 941 43638 3275
rect 49435 3348 49566 3405
rect 43572 939 44012 941
rect 43572 875 44027 939
rect 43870 0 44027 875
rect 49435 849 49492 3348
rect 50117 3323 50175 3519
rect 49906 3267 50175 3323
rect 50648 3328 50713 3522
rect 50648 3271 50917 3328
rect 49906 849 49962 3267
rect 50299 2937 50305 2977
rect 50860 2937 50917 3271
rect 51266 3256 51332 3514
rect 57322 3279 57387 3555
rect 51266 3210 51468 3256
rect 51266 3190 51469 3210
rect 50859 1673 50916 2937
rect 50859 1612 50986 1673
rect 49376 0 49533 849
rect 49847 0 50004 849
rect 50126 0 50282 1202
rect 50641 0 50797 1200
rect 50929 849 50986 1612
rect 51405 849 51469 3190
rect 57174 3195 57387 3279
rect 57929 3281 57994 3521
rect 57929 3203 58397 3281
rect 57174 849 57240 3195
rect 50921 0 51077 849
rect 51392 0 51548 849
rect 57098 0 57255 849
rect 57686 0 57843 1199
rect 58240 1006 58397 3203
rect 58160 861 58397 1006
rect 59066 2825 59766 7458
rect 59066 2581 59767 2825
rect 58160 0 58317 861
rect 59066 197 59766 2581
<< metal3 >>
rect 1018 44560 1717 44986
rect 1874 44560 2574 44986
rect 2896 44560 3595 44986
rect 3752 44560 4452 44986
rect 4926 44560 5625 44986
rect 5782 44560 6482 44986
rect 6676 44560 7375 44986
rect 7532 44560 8232 44986
rect 8834 44560 9533 44986
rect 9690 44560 10390 44986
rect 10456 44560 11155 44986
rect 11312 44560 12012 44986
rect 12742 44560 13441 44986
rect 13598 44560 14298 44986
rect 14457 44560 15156 44986
rect 16080 44560 16780 44986
rect 16937 44560 17636 44986
rect 17761 44560 18461 44986
rect 18600 44560 19299 44986
rect 19664 44560 20364 44986
rect 20641 44560 21341 44986
rect 21497 44560 22196 44986
rect 22817 44560 23517 44986
rect 23967 44560 24667 44986
rect 24790 44560 25489 44986
rect 26014 44560 26714 44986
rect 27009 44560 27708 44986
rect 28068 44560 28768 44986
rect 28861 44560 29560 44986
rect 29851 44560 30551 44986
rect 30749 44560 31449 44986
rect 31548 44560 32247 44986
rect 32419 44560 33118 44986
rect 33275 44560 33975 44986
rect 34231 44560 34930 44986
rect 35476 44560 36176 44986
rect 36798 44560 37497 44986
rect 37983 44560 38682 44986
rect 39343 44560 40043 44986
rect 40283 44663 40982 44986
rect 41104 44663 41804 44986
rect 42104 44560 42803 44986
rect 42960 44560 43660 44986
rect 44399 44560 45098 44986
rect 45255 44560 45955 44986
rect 46012 44560 46711 44986
rect 46868 44560 47568 44986
rect 48179 44560 48878 44986
rect 49035 44560 49735 44986
rect 49920 44560 50619 44986
rect 50776 44560 51476 44986
rect 51959 44560 52658 44986
rect 52815 44560 53515 44986
rect 53828 44560 54527 44986
rect 54684 44560 55384 44986
rect 55860 44560 56559 44986
rect 57166 44560 57866 44986
rect 58023 44560 58722 44986
rect 59066 44560 59765 44986
rect 42104 44559 42612 44560
rect 0 43726 60260 44426
rect 0 43160 709 43650
rect 19042 43335 19445 43476
rect 37782 43311 41389 43452
rect 0 42530 709 43020
rect 38000 43018 42103 43159
rect 59550 43137 60260 43626
rect 59550 42547 60260 43037
rect 0 41948 709 42438
rect 59550 41945 60260 42435
rect 0 41318 709 41808
rect 59550 41335 60260 41825
rect 0 40736 709 41226
rect 59550 40733 60260 41223
rect 0 40106 709 40596
rect 59550 40123 60260 40613
rect 0 39524 709 40014
rect 59550 39521 60260 40011
rect 0 38894 709 39384
rect 59550 38911 60260 39401
rect 0 38312 709 38802
rect 59550 38309 60260 38799
rect 0 37682 709 38172
rect 59550 37699 60260 38189
rect 0 37100 709 37590
rect 59550 37097 60260 37587
rect 0 36470 709 36960
rect 59550 36487 60260 36977
rect 0 35888 709 36378
rect 59550 35885 60260 36375
rect 0 35258 709 35748
rect 59550 35275 60260 35765
rect 0 34676 709 35166
rect 59550 34673 60260 35163
rect 0 34046 709 34536
rect 59550 34063 60260 34553
rect 0 33464 709 33929
rect 59550 33461 60260 33951
rect 0 32834 709 33324
rect 59550 32851 60260 33341
rect 0 32252 709 32742
rect 59550 32249 60260 32739
rect 0 31622 709 32112
rect 59550 31639 60260 32129
rect 0 31040 709 31530
rect 59550 31037 60260 31527
rect 0 30410 709 30900
rect 59550 30427 60260 30917
rect 0 29828 709 30318
rect 59550 29825 60260 30315
rect 0 29198 709 29688
rect 59550 29215 60260 29705
rect 0 28616 709 29106
rect 59550 28613 60260 29103
rect 0 27986 709 28476
rect 59550 28003 60260 28493
rect 0 27404 709 27894
rect 59550 27401 60260 27891
rect 0 26774 709 27264
rect 59550 26791 60260 27281
rect 0 26192 709 26682
rect 59550 26189 60260 26679
rect 0 25562 709 26052
rect 59550 25579 60260 26069
rect 0 24980 709 25470
rect 59551 25438 60260 25467
rect 59550 24977 60260 25438
rect 0 24350 709 24840
rect 59550 24367 60260 24857
rect 0 23768 709 24258
rect 59551 24216 60260 24255
rect 59550 23765 60260 24216
rect 0 23138 709 23628
rect 0 22270 709 22823
rect 17459 22404 19481 22606
rect 17529 22270 19481 22404
rect 0 19036 709 21982
rect 17529 20845 19049 21981
rect 25804 21843 26420 23239
rect 59550 23155 60260 23645
rect 40953 22270 42191 22606
rect 59550 22270 60260 22872
rect 19170 20900 20250 21479
rect 39294 20899 40415 21479
rect 40535 20764 42798 21981
rect 18740 20634 20249 20764
rect 39294 20715 42798 20764
rect 18740 20296 20250 20634
rect 39294 20303 40845 20715
rect 17977 19659 20267 20240
rect 39328 19663 41466 20241
rect 18740 19234 20247 19578
rect 39335 19234 40845 19567
rect 16863 19051 20250 19234
rect 16863 19036 20252 19051
rect 18740 18828 20252 19036
rect 39335 19036 42942 19234
rect 59550 19036 60260 21982
rect 0 17379 709 18766
rect 17186 17708 18529 18769
rect 18740 18083 20250 18828
rect 39335 18086 40845 19036
rect 17186 17388 19479 17708
rect 40949 17695 43331 18760
rect 40106 17376 43331 17695
rect 59550 17379 60260 18766
rect 16965 17105 18683 17255
rect 16965 16869 18466 17020
rect 16965 16626 18289 16776
rect 16965 16385 18118 16536
rect 19167 16486 20789 16963
rect 40531 16407 40852 16410
rect 16963 16157 17940 16307
rect 16963 15912 17771 16062
rect 18739 16038 40853 16407
rect 0 14971 709 15671
rect 16963 15667 17606 15817
rect 16973 15421 17411 15572
rect 18739 15281 19046 16038
rect 16825 14972 19046 15281
rect 19172 15504 40417 15965
rect 16825 14971 18720 14972
rect 19172 14754 19482 15504
rect 40102 14858 40417 15504
rect 19170 14730 19482 14754
rect 16862 14572 19482 14730
rect 0 13871 711 14571
rect 16825 14418 19482 14572
rect 40103 14702 40417 14858
rect 40531 15281 40852 16038
rect 40531 14856 43362 15281
rect 59550 14971 60260 15671
rect 16825 14253 17418 14418
rect 40103 14388 42858 14702
rect 17533 13771 42273 14310
rect 42402 14255 42858 14388
rect 59551 14172 60260 14572
rect 59550 13871 60260 14172
rect 17533 13552 18072 13771
rect 0 11642 709 13537
rect 16825 13013 18072 13552
rect 18538 13446 20582 13606
rect 39004 13445 41081 13605
rect 41734 13555 42273 13771
rect 18345 13208 20582 13368
rect 39004 13207 41321 13367
rect 18174 12970 20582 13130
rect 39004 12969 41528 13129
rect 41734 13016 42729 13555
rect 18001 12732 20582 12892
rect 39004 12731 41738 12891
rect 17821 12494 20582 12654
rect 39004 12493 41945 12653
rect 17642 12256 20582 12416
rect 39004 12255 42166 12415
rect 17483 12018 20582 12178
rect 39004 12017 42360 12177
rect 17282 11780 20582 11940
rect 39004 11779 42576 11939
rect 59550 11642 60260 13550
rect 0 9590 709 11442
rect 38898 11343 42993 11446
rect 16877 9947 19479 11184
rect 38898 10274 42994 11343
rect 16877 9635 20636 9947
rect 0 8025 709 9465
rect 16832 8848 19049 9530
rect 19170 9066 20636 9635
rect 40098 9585 42733 10274
rect 42991 9969 42994 10274
rect 59550 9591 60260 11442
rect 38824 9461 39860 9501
rect 38824 9177 43638 9461
rect 16832 8041 20637 8848
rect 38824 8807 40914 9177
rect 38824 8239 43638 8807
rect 16832 8037 18587 8041
rect 38824 7982 40880 8239
rect 59550 8002 60260 9462
rect 0 6723 709 7645
rect 16832 6728 19479 7650
rect 38902 7648 40882 7840
rect 38902 7313 43594 7648
rect 36220 6909 39257 6971
rect 36220 6652 36282 6909
rect 39195 6626 39257 6909
rect 40106 6728 43594 7313
rect 59550 6724 60260 7646
rect 2933 6564 20454 6626
rect 39195 6564 43501 6626
rect 20393 6336 20454 6564
rect 40415 6381 43594 6448
rect 20393 6274 29159 6336
rect 0 5306 709 6260
rect 16832 5312 20110 6266
rect 29097 6089 29159 6274
rect 29097 6027 35046 6089
rect 38832 6034 40415 6244
rect 18434 5311 20110 5312
rect 0 3963 709 5093
rect 16541 4922 19479 5093
rect 16537 4729 19479 4922
rect 19635 5060 20110 5311
rect 38836 5092 40415 6034
rect 40536 5522 43594 6264
rect 40536 5311 42899 5522
rect 59550 5305 60260 6259
rect 38836 5078 43922 5092
rect 19635 4858 20696 5060
rect 38833 4881 43922 5078
rect 19727 4668 20272 4751
rect 16537 4572 20273 4668
rect 16541 4497 20273 4572
rect 16537 4330 20273 4497
rect 39245 4653 39871 4792
rect 40105 4730 43922 4881
rect 19727 4324 20272 4330
rect 39245 4325 43922 4653
rect 16537 4019 16541 4190
rect 16580 3962 20911 4265
rect 38836 3958 43700 4261
rect 59550 3962 60260 5092
rect 0 2844 709 3870
rect 16580 3548 19049 3867
rect 40536 3606 43699 3867
rect 40536 3545 43700 3606
rect 40538 3102 43081 3242
rect 40538 2984 43702 3102
rect 42823 2844 43702 2984
rect 59550 2841 60260 3870
rect 40097 2645 42575 2785
rect 0 1994 709 2637
rect 40097 2527 43700 2645
rect 42324 2387 43700 2527
rect 17006 2083 43067 2144
rect 59570 1995 60260 2639
rect 58724 1994 60260 1995
rect 0 1750 60260 1994
rect 0 1749 59613 1750
rect 0 1748 58724 1749
rect 50835 1709 50913 1748
rect 40536 1562 43700 1567
rect 58724 1562 58933 1563
rect 0 862 60260 1562
rect 493 818 1194 862
rect 494 0 1194 818
rect 1427 0 2127 862
rect 2409 0 3109 862
rect 3249 0 3949 311
rect 4089 0 4789 862
rect 4929 0 5629 862
rect 5769 0 6469 862
rect 6609 0 7309 311
rect 7449 0 8149 862
rect 8710 0 9410 862
rect 9969 0 10669 862
rect 10809 0 11509 311
rect 11649 0 12349 862
rect 12489 0 13189 862
rect 13329 0 14029 862
rect 14169 0 14869 311
rect 15337 0 16037 862
rect 16177 0 16877 862
rect 17087 0 17787 862
rect 17997 0 18697 862
rect 18907 0 19607 862
rect 19817 0 20517 862
rect 20727 0 21427 862
rect 21926 0 22626 311
rect 23115 0 23815 311
rect 24381 0 25081 311
rect 25221 0 25921 862
rect 26619 0 27319 311
rect 27459 0 28159 862
rect 28863 0 29563 311
rect 29703 0 30403 862
rect 30543 0 31243 311
rect 31383 0 32083 862
rect 32223 0 32923 311
rect 33063 0 33763 862
rect 33996 0 34696 862
rect 34913 0 35613 862
rect 35863 0 36563 311
rect 38120 0 38820 862
rect 39030 0 39730 862
rect 39940 841 44306 862
rect 39940 0 40640 841
rect 40850 0 41550 841
rect 41760 0 42460 841
rect 42670 0 43370 841
rect 43606 0 44306 841
rect 44752 0 45452 311
rect 45592 0 46292 862
rect 46432 0 47132 862
rect 47272 0 47972 862
rect 48112 0 48812 311
rect 48952 0 49652 862
rect 50211 0 50911 862
rect 51472 0 52172 862
rect 52312 0 53012 311
rect 53152 0 53852 862
rect 53992 0 54692 862
rect 54832 0 55532 862
rect 55672 0 56372 311
rect 56712 0 57412 862
rect 57693 0 58393 862
rect 59066 0 59766 862
use 3v256x8M8W_PWR_3v256x8m81  3v256x8M8W_PWR_3v256x8m81_0
timestamp 1765833452
transform 1 0 0 0 1 -1905
box 1338 9885 58383 24803
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_0
timestamp 1765475971
transform 0 1 1382 -1 0 1003
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_1
timestamp 1765475971
transform 0 1 2094 -1 0 1003
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_2
timestamp 1765475971
transform 0 1 8674 -1 0 1003
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_3
timestamp 1765475971
transform 0 1 8918 -1 0 1003
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_4
timestamp 1765475971
transform 0 1 9218 -1 0 1003
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_5
timestamp 1765475971
transform 0 1 9542 -1 0 1003
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_6
timestamp 1765475971
transform 0 1 16454 -1 0 1003
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_7
timestamp 1765475971
transform 0 1 17173 -1 0 1003
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_8
timestamp 1765475971
transform 0 1 19647 -1 0 1451
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_9
timestamp 1765475971
transform 0 1 43361 -1 0 1002
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_10
timestamp 1765475971
transform 0 1 49940 -1 0 1002
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_11
timestamp 1765475971
transform 0 1 50240 -1 0 1002
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_12
timestamp 1765475971
transform 0 1 50676 -1 0 1002
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_13
timestamp 1765475971
transform 0 1 50976 -1 0 1002
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_14
timestamp 1765475971
transform 0 1 57766 -1 0 1002
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_15
timestamp 1765475971
transform 0 1 42488 -1 0 1002
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_16
timestamp 1765475971
transform 0 1 35315 -1 0 1504
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_17
timestamp 1765475971
transform 0 1 28489 -1 0 1461
box -53 -92 53 93
use antenna_tiedown_3v256x8m81  antenna_tiedown_3v256x8m81_18
timestamp 1765475971
transform 0 1 58317 -1 0 1002
box -53 -92 53 93
use control_3v256x8_3v256x8m81  control_3v256x8_3v256x8m81_0
timestamp 1765847097
transform 1 0 19273 0 1 1392
box -2537 648 22252 21087
use G_ring_3v256x8m81  G_ring_3v256x8m81_0
timestamp 1763766357
transform 1 0 197 0 1 -1905
box 0 1905 59871 46326
use GF018_3v256x8M8WM1_lef_3v256x8m81  GF018_3v256x8M8WM1_lef_3v256x8m81_0
timestamp 1764698730
transform 1 0 0 0 1 0
box 0 0 60260 44986
use lcol4_256_3v256x8m81  lcol4_256_3v256x8m81_0
timestamp 1765899468
transform 1 0 2044 0 1 1608
box -830 -478 15967 41903
use M1_PSUB4310591302010_3v256x8m81  M1_PSUB4310591302010_3v256x8m81_0
timestamp 1763766357
transform 1 0 37597 0 1 2041
box -2018 -800 2018 800
use M1_PSUB4310591302014_3v256x8m81  M1_PSUB4310591302014_3v256x8m81_0
timestamp 1763766357
transform 1 0 24082 0 1 2041
box -4048 -800 4048 800
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_0
timestamp 1763766357
transform 1 0 39671 0 1 24000
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_1
timestamp 1763766357
transform 1 0 39671 0 1 25212
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_2
timestamp 1763766357
transform 1 0 39671 0 1 26425
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_3
timestamp 1763766357
transform 1 0 39671 0 1 27636
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_4
timestamp 1763766357
transform 1 0 39671 0 1 28848
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_5
timestamp 1763766357
transform 1 0 39671 0 1 30060
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_6
timestamp 1763766357
transform 1 0 39671 0 1 31272
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_7
timestamp 1763766357
transform 1 0 19914 0 1 31273
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_8
timestamp 1763766357
transform 1 0 19914 0 1 30060
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_9
timestamp 1763766357
transform 1 0 19914 0 1 28848
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_10
timestamp 1763766357
transform 1 0 19914 0 1 27636
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_11
timestamp 1763766357
transform 1 0 19914 0 1 24003
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_12
timestamp 1763766357
transform 1 0 19914 0 1 25213
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_13
timestamp 1763766357
transform 1 0 19914 0 1 26423
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_29
timestamp 1763766357
transform 1 0 19914 0 1 43392
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_30
timestamp 1763766357
transform 1 0 19914 0 1 42180
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_31
timestamp 1763766357
transform 1 0 19914 0 1 40968
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_32
timestamp 1763766357
transform 1 0 19914 0 1 39756
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_33
timestamp 1763766357
transform 1 0 19914 0 1 38544
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_34
timestamp 1763766357
transform 1 0 19914 0 1 37332
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_35
timestamp 1763766357
transform 1 0 19914 0 1 36120
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_36
timestamp 1763766357
transform 1 0 19914 0 1 34908
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_37
timestamp 1763766357
transform 1 0 19914 0 1 33696
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_38
timestamp 1763766357
transform 1 0 19914 0 1 32484
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_39
timestamp 1763766357
transform 1 0 19914 0 1 43392
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_45
timestamp 1763766357
transform 1 0 39671 0 1 32484
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_46
timestamp 1763766357
transform 1 0 39671 0 1 33696
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_47
timestamp 1763766357
transform 1 0 39671 0 1 34908
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_48
timestamp 1763766357
transform 1 0 39671 0 1 36120
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_49
timestamp 1763766357
transform 1 0 39671 0 1 37332
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_50
timestamp 1763766357
transform 1 0 39671 0 1 38544
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_51
timestamp 1763766357
transform 1 0 39671 0 1 39756
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_52
timestamp 1763766357
transform 1 0 39671 0 1 40968
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_53
timestamp 1763766357
transform 1 0 39671 0 1 42180
box -487 -46 487 46
use M2_M1$$199747628_3v256x8m81  M2_M1$$199747628_3v256x8m81_54
timestamp 1763766357
transform 1 0 39671 0 1 43392
box -487 -46 487 46
use M2_M1$$201260076_3v256x8m81  M2_M1$$201260076_3v256x8m81_0
timestamp 1763766357
transform -1 0 40260 0 1 11653
box -119 -9872 119 9872
use M2_M1$$201260076_3v256x8m81  M2_M1$$201260076_3v256x8m81_1
timestamp 1763766357
transform -1 0 40691 0 1 11653
box -119 -9872 119 9872
use M2_M1$$201260076_3v256x8m81  M2_M1$$201260076_3v256x8m81_2
timestamp 1763766357
transform 1 0 19325 0 1 11653
box -119 -9872 119 9872
use M2_M1$$201260076_3v256x8m81  M2_M1$$201260076_3v256x8m81_3
timestamp 1763766357
transform 1 0 18895 0 1 11653
box -119 -9872 119 9872
use M2_M1431059130200_3v256x8m81  M2_M1431059130200_3v256x8m81_0
timestamp 1765833244
transform 1 0 43359 0 1 1154
box -63 -34 63 34
use M2_M1431059130200_3v256x8m81  M2_M1431059130200_3v256x8m81_1
timestamp 1765833244
transform 1 0 34990 0 1 4221
box -63 -34 63 34
use M2_M1431059130200_3v256x8m81  M2_M1431059130200_3v256x8m81_2
timestamp 1765833244
transform 1 0 57765 0 1 1164
box -63 -34 63 34
use M2_M1431059130200_3v256x8m81  M2_M1431059130200_3v256x8m81_3
timestamp 1765833244
transform 1 0 36212 0 1 3416
box -63 -34 63 34
use M2_M1431059130200_3v256x8m81  M2_M1431059130200_3v256x8m81_4
timestamp 1765833244
transform 1 0 50720 0 1 1163
box -63 -34 63 34
use M2_M1431059130200_3v256x8m81  M2_M1431059130200_3v256x8m81_5
timestamp 1765833244
transform 1 0 50205 0 1 1163
box -63 -34 63 34
use M2_M1431059130200_3v256x8m81  M2_M1431059130200_3v256x8m81_6
timestamp 1765833244
transform 1 0 16461 0 1 1164
box -63 -34 63 34
use M2_M1431059130200_3v256x8m81  M2_M1431059130200_3v256x8m81_7
timestamp 1765833244
transform 1 0 9246 0 1 1164
box -63 -34 63 34
use M2_M1431059130200_3v256x8m81  M2_M1431059130200_3v256x8m81_8
timestamp 1765833244
transform 1 0 8901 0 1 1164
box -63 -34 63 34
use M2_M1431059130200_3v256x8m81  M2_M1431059130200_3v256x8m81_9
timestamp 1765833244
transform 1 0 2106 0 1 1163
box -63 -34 63 34
use M2_M1431059130200_3v256x8m81  M2_M1431059130200_3v256x8m81_10
timestamp 1765833244
transform 1 0 28490 0 1 2038
box -63 -34 63 34
use M2_M1431059130203_3v256x8m81  M2_M1431059130203_3v256x8m81_0
timestamp 1763766357
transform 1 0 18271 0 1 22438
box -200 -156 200 156
use M2_M1431059130204_3v256x8m81  M2_M1431059130204_3v256x8m81_0
timestamp 1763766357
transform 1 0 18293 0 1 43409
box -200 -113 200 113
use M2_M1431059130204_3v256x8m81  M2_M1431059130204_3v256x8m81_1
timestamp 1763766357
transform 1 0 41198 0 1 43479
box -200 -113 200 113
use M2_M1431059130208_3v256x8m81  M2_M1431059130208_3v256x8m81_0
timestamp 1765833244
transform 1 0 41860 0 1 22892
box -34 -63 34 63
use M2_M14310591302012_3v256x8m81  M2_M14310591302012_3v256x8m81_0
timestamp 1763766357
transform 1 0 19319 0 1 22439
box -113 -156 113 156
use M2_M14310591302012_3v256x8m81  M2_M14310591302012_3v256x8m81_1
timestamp 1763766357
transform 1 0 20383 0 1 1116
box -113 -156 113 156
use m2m3_3v256x8m81  m2m3_3v256x8m81_0
timestamp 1763766357
transform 1 0 41027 0 1 10080
box -75 1710 1856 7189
use M3_M2$$201248812_3v256x8m81  M3_M2$$201248812_3v256x8m81_0
timestamp 1763766357
transform -1 0 40691 0 1 8723
box -119 -732 119 732
use M3_M2$$201248812_3v256x8m81  M3_M2$$201248812_3v256x8m81_1
timestamp 1763766357
transform -1 0 40260 0 1 10464
box -119 -732 119 732
use M3_M2$$201248812_3v256x8m81  M3_M2$$201248812_3v256x8m81_2
timestamp 1763766357
transform 1 0 19325 0 1 10429
box -119 -732 119 732
use M3_M2$$201248812_3v256x8m81  M3_M2$$201248812_3v256x8m81_3
timestamp 1763766357
transform 1 0 18895 0 1 8783
box -119 -732 119 732
use M3_M2$$201249836_3v256x8m81  M3_M2$$201249836_3v256x8m81_0
timestamp 1763766357
transform -1 0 40260 0 1 7368
box -119 -427 119 427
use M3_M2$$201249836_3v256x8m81  M3_M2$$201249836_3v256x8m81_1
timestamp 1763766357
transform -1 0 40691 0 1 5799
box -119 -427 119 427
use M3_M2$$201249836_3v256x8m81  M3_M2$$201249836_3v256x8m81_2
timestamp 1763766357
transform 1 0 19325 0 1 7188
box -119 -427 119 427
use M3_M2$$201249836_3v256x8m81  M3_M2$$201249836_3v256x8m81_3
timestamp 1763766357
transform 1 0 18895 0 1 5819
box -119 -427 119 427
use M3_M2$$201250860_3v256x8m81  M3_M2$$201250860_3v256x8m81_0
timestamp 1763766357
transform -1 0 39553 0 1 4548
box -266 -198 266 198
use M3_M2$$201250860_3v256x8m81  M3_M2$$201250860_3v256x8m81_1
timestamp 1763766357
transform 1 0 20002 0 1 4539
box -266 -198 266 198
use M3_M2$$201251884_3v256x8m81  M3_M2$$201251884_3v256x8m81_0
timestamp 1763766357
transform 1 0 26112 0 1 23192
box -266 -46 266 46
use M3_M2$$201252908_3v256x8m81  M3_M2$$201252908_3v256x8m81_0
timestamp 1765833244
transform 1 0 20180 0 1 2659
box -45 -122 45 123
use M3_M2$$201253932_3v256x8m81  M3_M2$$201253932_3v256x8m81_0
timestamp 1763766357
transform 1 0 40260 0 1 5708
box -119 -808 119 511
use M3_M2$$201254956_3v256x8m81  M3_M2$$201254956_3v256x8m81_0
timestamp 1763766357
transform 1 0 19325 0 1 9242
box -119 -151 119 351
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_0
timestamp 1763766357
transform 1 0 19914 0 1 32484
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_1
timestamp 1763766357
transform 1 0 39671 0 1 25212
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_2
timestamp 1763766357
transform 1 0 39671 0 1 26425
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_3
timestamp 1763766357
transform 1 0 39671 0 1 27636
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_4
timestamp 1763766357
transform 1 0 39671 0 1 28848
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_5
timestamp 1763766357
transform 1 0 39671 0 1 30060
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_6
timestamp 1763766357
transform 1 0 39671 0 1 31272
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_7
timestamp 1763766357
transform 1 0 19914 0 1 31272
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_8
timestamp 1763766357
transform 1 0 19914 0 1 30060
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_9
timestamp 1763766357
transform 1 0 19914 0 1 28848
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_10
timestamp 1763766357
transform 1 0 19914 0 1 27636
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_11
timestamp 1763766357
transform 1 0 19914 0 1 26423
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_12
timestamp 1763766357
transform 1 0 19914 0 1 25215
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_13
timestamp 1763766357
transform 1 0 19914 0 1 24003
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_23
timestamp 1763766357
transform 1 0 19914 0 1 43392
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_24
timestamp 1763766357
transform 1 0 19914 0 1 42180
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_25
timestamp 1763766357
transform 1 0 19914 0 1 40968
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_26
timestamp 1763766357
transform 1 0 19914 0 1 39756
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_27
timestamp 1763766357
transform 1 0 19914 0 1 38544
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_28
timestamp 1763766357
transform 1 0 19914 0 1 37332
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_29
timestamp 1763766357
transform 1 0 19914 0 1 36120
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_30
timestamp 1763766357
transform 1 0 19914 0 1 34908
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_31
timestamp 1763766357
transform 1 0 19914 0 1 33696
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_32
timestamp 1763766357
transform 1 0 19914 0 1 32484
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_33
timestamp 1763766357
transform 1 0 19914 0 1 43392
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_40
timestamp 1763766357
transform 1 0 39671 0 1 32484
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_41
timestamp 1763766357
transform 1 0 39671 0 1 33696
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_42
timestamp 1763766357
transform 1 0 39671 0 1 34908
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_43
timestamp 1763766357
transform 1 0 39671 0 1 36120
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_44
timestamp 1763766357
transform 1 0 39671 0 1 37332
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_45
timestamp 1763766357
transform 1 0 39671 0 1 38544
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_46
timestamp 1763766357
transform 1 0 39671 0 1 39756
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_47
timestamp 1763766357
transform 1 0 39671 0 1 40968
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_48
timestamp 1763766357
transform 1 0 39671 0 1 42180
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_65
timestamp 1763766357
transform 1 0 39671 0 1 43390
box -487 -46 487 46
use M3_M2$$201258028_3v256x8m81  M3_M2$$201258028_3v256x8m81_66
timestamp 1763766357
transform 1 0 39671 0 1 24000
box -487 -46 487 46
use M3_M2$$201412652_3v256x8m81  M3_M2$$201412652_3v256x8m81_0
timestamp 1763766357
transform -1 0 40260 0 1 19942
box -119 -275 119 275
use M3_M2$$201412652_3v256x8m81  M3_M2$$201412652_3v256x8m81_1
timestamp 1763766357
transform -1 0 40260 0 1 21185
box -119 -275 119 275
use M3_M2$$201412652_3v256x8m81  M3_M2$$201412652_3v256x8m81_2
timestamp 1763766357
transform 1 0 19325 0 1 21185
box -119 -275 119 275
use M3_M2$$201412652_3v256x8m81  M3_M2$$201412652_3v256x8m81_3
timestamp 1763766357
transform 1 0 19325 0 1 19921
box -119 -275 119 275
use M3_M2$$201413676_3v256x8m81  M3_M2$$201413676_3v256x8m81_0
timestamp 1763766357
transform -1 0 40691 0 1 20504
box -119 -158 119 198
use M3_M2$$201413676_3v256x8m81  M3_M2$$201413676_3v256x8m81_1
timestamp 1763766357
transform 1 0 18895 0 1 20514
box -119 -158 119 198
use M3_M2$$201413676_3v256x8m81  M3_M2$$201413676_3v256x8m81_2
timestamp 1763766357
transform 1 0 19325 0 1 4888
box -119 -158 119 198
use M3_M2$$201414700_3v256x8m81  M3_M2$$201414700_3v256x8m81_0
timestamp 1763766357
transform -1 0 40691 0 1 21349
box -119 -479 119 579
use M3_M2$$201414700_3v256x8m81  M3_M2$$201414700_3v256x8m81_1
timestamp 1763766357
transform 1 0 18895 0 1 21349
box -119 -479 119 579
use M3_M2$$201415724_3v256x8m81  M3_M2$$201415724_3v256x8m81_0
timestamp 1763766357
transform -1 0 40691 0 1 18675
box -119 -584 119 884
use M3_M2$$201415724_3v256x8m81  M3_M2$$201415724_3v256x8m81_1
timestamp 1763766357
transform 1 0 18895 0 1 18679
box -119 -584 119 884
use M3_M2$$201416748_3v256x8m81  M3_M2$$201416748_3v256x8m81_0
timestamp 1765833244
transform -1 0 40260 0 1 2655
box -119 -123 119 123
use M3_M2$$201416748_3v256x8m81  M3_M2$$201416748_3v256x8m81_1
timestamp 1765833244
transform -1 0 40691 0 1 3716
box -119 -123 119 123
use M3_M2$$201416748_3v256x8m81  M3_M2$$201416748_3v256x8m81_2
timestamp 1765833244
transform -1 0 40260 0 1 4123
box -119 -123 119 123
use M3_M2$$201416748_3v256x8m81  M3_M2$$201416748_3v256x8m81_3
timestamp 1765833244
transform -1 0 40691 0 1 3113
box -119 -123 119 123
use M3_M2$$201416748_3v256x8m81  M3_M2$$201416748_3v256x8m81_4
timestamp 1765833244
transform -1 0 40260 0 1 17535
box -119 -123 119 123
use M3_M2$$201416748_3v256x8m81  M3_M2$$201416748_3v256x8m81_5
timestamp 1765833244
transform 1 0 19325 0 1 2660
box -119 -123 119 123
use M3_M2$$201416748_3v256x8m81  M3_M2$$201416748_3v256x8m81_6
timestamp 1765833244
transform 1 0 18895 0 1 3143
box -119 -123 119 123
use M3_M2$$201416748_3v256x8m81  M3_M2$$201416748_3v256x8m81_7
timestamp 1765833244
transform 1 0 19325 0 1 4114
box -119 -123 119 123
use M3_M2$$201416748_3v256x8m81  M3_M2$$201416748_3v256x8m81_8
timestamp 1765833244
transform 1 0 18895 0 1 3707
box -119 -123 119 123
use M3_M2$$201416748_3v256x8m81  M3_M2$$201416748_3v256x8m81_9
timestamp 1765833244
transform 1 0 19325 0 1 17548
box -119 -123 119 123
use M3_M2$$201416748_3v256x8m81  M3_M2$$201416748_3v256x8m81_10
timestamp 1765833244
transform 1 0 19325 0 1 16741
box -119 -123 119 123
use M3_M2$$204143660_3v256x8m81  M3_M2$$204143660_3v256x8m81_0
timestamp 1763766357
transform 1 0 29305 0 1 42786
box -45 -46 171 46
use M3_M2431059130201_3v256x8m81  M3_M2431059130201_3v256x8m81_0
timestamp 1765833244
transform 0 -1 34983 1 0 6042
box -35 -63 35 63
use M3_M2431059130201_3v256x8m81  M3_M2431059130201_3v256x8m81_1
timestamp 1765833244
transform 1 0 36255 0 1 6718
box -35 -63 35 63
use M3_M2431059130202_3v256x8m81  M3_M2431059130202_3v256x8m81_0
timestamp 1763766357
transform 1 0 18271 0 1 22439
box -200 -156 200 156
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_0
timestamp 1763766357
transform 1 0 40689 0 1 14158
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_1
timestamp 1763766357
transform 1 0 40689 0 1 13917
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_2
timestamp 1763766357
transform 1 0 17352 0 1 11860
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_3
timestamp 1763766357
transform 1 0 17527 0 1 15741
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_4
timestamp 1763766357
transform 1 0 17546 0 1 12098
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_5
timestamp 1763766357
transform 1 0 17696 0 1 15986
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_6
timestamp 1763766357
transform 1 0 17715 0 1 12322
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_7
timestamp 1763766357
transform 1 0 17872 0 1 16230
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_8
timestamp 1763766357
transform 1 0 17891 0 1 12584
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_9
timestamp 1763766357
transform 1 0 18050 0 1 16462
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_10
timestamp 1763766357
transform 1 0 18069 0 1 12817
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_11
timestamp 1763766357
transform 1 0 18225 0 1 16696
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_12
timestamp 1763766357
transform 1 0 18245 0 1 13057
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_13
timestamp 1763766357
transform 1 0 18400 0 1 16939
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_14
timestamp 1763766357
transform 1 0 18420 0 1 13281
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_15
timestamp 1763766357
transform 1 0 18611 0 1 17173
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_16
timestamp 1763766357
transform 1 0 18611 0 1 13523
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_17
timestamp 1763766357
transform 1 0 18902 0 1 14168
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_18
timestamp 1763766357
transform 1 0 18902 0 1 13927
box -63 -63 63 63
use M3_M2431059130205_3v256x8m81  M3_M2431059130205_3v256x8m81_19
timestamp 1763766357
transform 1 0 17335 0 1 15496
box -63 -63 63 63
use M3_M2431059130206_3v256x8m81  M3_M2431059130206_3v256x8m81_0
timestamp 1763766357
transform 1 0 19319 0 1 22439
box -113 -156 113 156
use M3_M2431059130207_3v256x8m81  M3_M2431059130207_3v256x8m81_0
timestamp 1765833244
transform 1 0 30716 0 1 2114
box -63 -35 63 35
use M3_M2431059130209_3v256x8m81  M3_M2431059130209_3v256x8m81_0
timestamp 1763766357
transform 1 0 41204 0 1 20097
box -200 -113 200 113
use M3_M2431059130209_3v256x8m81  M3_M2431059130209_3v256x8m81_1
timestamp 1763766357
transform 1 0 41204 0 1 19825
box -200 -113 200 113
use M3_M2431059130209_3v256x8m81  M3_M2431059130209_3v256x8m81_2
timestamp 1763766357
transform 1 0 18271 0 1 20101
box -200 -113 200 113
use M3_M2431059130209_3v256x8m81  M3_M2431059130209_3v256x8m81_3
timestamp 1763766357
transform 1 0 18271 0 1 19782
box -200 -113 200 113
use M3_M2431059130209_3v256x8m81  M3_M2431059130209_3v256x8m81_4
timestamp 1763766357
transform 1 0 18293 0 1 43409
box -200 -113 200 113
use M3_M2431059130209_3v256x8m81  M3_M2431059130209_3v256x8m81_5
timestamp 1763766357
transform 1 0 41198 0 1 43479
box -200 -113 200 113
use M3_M24310591302011_3v256x8m81  M3_M24310591302011_3v256x8m81_0
timestamp 1763766357
transform 1 0 41207 0 1 22439
box -243 -156 243 156
use M3_M24310591302013_3v256x8m81  M3_M24310591302013_3v256x8m81_0
timestamp 1763766357
transform 1 0 40688 0 1 16046
box -99 -317 99 317
use M3_M24310591302013_3v256x8m81  M3_M24310591302013_3v256x8m81_1
timestamp 1763766357
transform 1 0 40246 0 1 15250
box -99 -317 99 317
use M3_M24310591302013_3v256x8m81  M3_M24310591302013_3v256x8m81_2
timestamp 1763766357
transform 1 0 18893 0 1 15456
box -99 -317 99 317
use M3_M24310591302013_3v256x8m81  M3_M24310591302013_3v256x8m81_3
timestamp 1763766357
transform 1 0 19324 0 1 14817
box -99 -317 99 317
use M3_M24310591302015_3v256x8m81  M3_M24310591302015_3v256x8m81_0
timestamp 1763766357
transform 1 0 41194 0 1 18104
box -200 -634 200 634
use M3_M24310591302015_3v256x8m81  M3_M24310591302015_3v256x8m81_1
timestamp 1763766357
transform 1 0 18276 0 1 18079
box -200 -634 200 634
use power_a_3v256x8m81  power_a_3v256x8m81_0
timestamp 1763766357
transform -1 0 48812 0 1 197
box 0 -197 700 700
use power_a_3v256x8m81  power_a_3v256x8m81_1
timestamp 1763766357
transform -1 0 56372 0 1 197
box 0 -197 700 700
use power_a_3v256x8m81  power_a_3v256x8m81_2
timestamp 1763766357
transform 1 0 52312 0 1 197
box 0 -197 700 700
use power_a_3v256x8m81  power_a_3v256x8m81_3
timestamp 1763766357
transform 1 0 32223 0 1 197
box 0 -197 700 700
use power_a_3v256x8m81  power_a_3v256x8m81_4
timestamp 1763766357
transform 1 0 36734 0 1 197
box 0 -197 700 700
use power_a_3v256x8m81  power_a_3v256x8m81_5
timestamp 1763766357
transform 1 0 30543 0 1 197
box 0 -197 700 700
use power_a_3v256x8m81  power_a_3v256x8m81_6
timestamp 1763766357
transform 1 0 35863 0 1 197
box 0 -197 700 700
use power_a_3v256x8m81  power_a_3v256x8m81_7
timestamp 1763766357
transform 1 0 44752 0 1 197
box 0 -197 700 700
use power_a_3v256x8m81  power_a_3v256x8m81_8
timestamp 1763766357
transform -1 0 23815 0 1 197
box 0 -197 700 700
use power_a_3v256x8m81  power_a_3v256x8m81_9
timestamp 1763766357
transform -1 0 22626 0 1 197
box 0 -197 700 700
use power_a_3v256x8m81  power_a_3v256x8m81_10
timestamp 1763766357
transform -1 0 7309 0 1 197
box 0 -197 700 700
use power_a_3v256x8m81  power_a_3v256x8m81_11
timestamp 1763766357
transform -1 0 14869 0 1 197
box 0 -197 700 700
use power_a_3v256x8m81  power_a_3v256x8m81_12
timestamp 1763766357
transform 1 0 28863 0 1 197
box 0 -197 700 700
use power_a_3v256x8m81  power_a_3v256x8m81_13
timestamp 1763766357
transform 1 0 10809 0 1 197
box 0 -197 700 700
use power_a_3v256x8m81  power_a_3v256x8m81_14
timestamp 1763766357
transform 1 0 24381 0 1 197
box 0 -197 700 700
use power_a_3v256x8m81  power_a_3v256x8m81_15
timestamp 1763766357
transform 1 0 3249 0 1 197
box 0 -197 700 700
use power_a_3v256x8m81  power_a_3v256x8m81_16
timestamp 1763766357
transform 1 0 26619 0 1 197
box 0 -197 700 700
use power_route_01_a_3v256x8m81  power_route_01_a_3v256x8m81_0
timestamp 1763766357
transform 1 0 10813 0 1 43285
box -357 441 1199 1701
use power_route_01_a_3v256x8m81  power_route_01_a_3v256x8m81_1
timestamp 1763766357
transform 1 0 7033 0 1 43285
box -357 441 1199 1701
use power_route_01_a_3v256x8m81  power_route_01_a_3v256x8m81_2
timestamp 1763766357
transform 1 0 3253 0 1 43285
box -357 441 1199 1701
use power_route_01_a_3v256x8m81  power_route_01_a_3v256x8m81_3
timestamp 1763766357
transform 1 0 52316 0 1 43285
box -357 441 1199 1701
use power_route_01_a_3v256x8m81  power_route_01_a_3v256x8m81_4
timestamp 1763766357
transform 1 0 48536 0 1 43285
box -357 441 1199 1701
use power_route_01_a_3v256x8m81  power_route_01_a_3v256x8m81_5
timestamp 1763766357
transform 1 0 44756 0 1 43285
box -357 441 1199 1701
use power_route_01_a_3v256x8m81  power_route_01_a_3v256x8m81_6
timestamp 1763766357
transform 1 0 32776 0 1 43285
box -357 441 1199 1701
use power_route_01_b_3v256x8m81  power_route_01_b_3v256x8m81_0
timestamp 1763766357
transform -1 0 29203 0 1 43285
box -357 441 342 1701
use power_route_01_b_3v256x8m81  power_route_01_b_3v256x8m81_1
timestamp 1763766357
transform -1 0 27351 0 1 43285
box -357 441 342 1701
use power_route_01_b_3v256x8m81  power_route_01_b_3v256x8m81_2
timestamp 1763766357
transform -1 0 25132 0 1 43285
box -357 441 342 1701
use power_route_01_b_3v256x8m81  power_route_01_b_3v256x8m81_3
timestamp 1763766357
transform -1 0 21839 0 1 43285
box -357 441 342 1701
use power_route_01_b_3v256x8m81  power_route_01_b_3v256x8m81_4
timestamp 1763766357
transform -1 0 18942 0 1 43285
box -357 441 342 1701
use power_route_01_b_3v256x8m81  power_route_01_b_3v256x8m81_5
timestamp 1763766357
transform -1 0 14799 0 1 43285
box -357 441 342 1701
use power_route_01_b_3v256x8m81  power_route_01_b_3v256x8m81_6
timestamp 1763766357
transform -1 0 56202 0 1 43285
box -357 441 342 1701
use power_route_01_b_3v256x8m81  power_route_01_b_3v256x8m81_7
timestamp 1763766357
transform -1 0 40625 0 1 43285
box -357 441 342 1701
use power_route_01_b_3v256x8m81  power_route_01_b_3v256x8m81_8
timestamp 1763766357
transform -1 0 59408 0 1 43285
box -357 441 342 1701
use power_route_01_b_3v256x8m81  power_route_01_b_3v256x8m81_9
timestamp 1763766357
transform -1 0 38325 0 1 43285
box -357 441 342 1701
use power_route_01_b_3v256x8m81  power_route_01_b_3v256x8m81_10
timestamp 1763766357
transform -1 0 34573 0 1 43285
box -357 441 342 1701
use power_route_01_b_3v256x8m81  power_route_01_b_3v256x8m81_11
timestamp 1763766357
transform -1 0 31890 0 1 43285
box -357 441 342 1701
use power_route_01_b_3v256x8m81  power_route_01_b_3v256x8m81_12
timestamp 1763766357
transform -1 0 37140 0 1 43285
box -357 441 342 1701
use power_route_01_c_3v256x8m81  power_route_01_c_3v256x8m81_0
timestamp 1763766357
transform -1 0 18810 0 1 43285
box 349 1275 1049 1701
use power_route_01_c_3v256x8m81  power_route_01_c_3v256x8m81_1
timestamp 1763766357
transform -1 0 29117 0 1 43285
box 349 1275 1049 1701
use power_route_01_c_3v256x8m81  power_route_01_c_3v256x8m81_2
timestamp 1763766357
transform -1 0 27063 0 1 43285
box 349 1275 1049 1701
use power_route_01_c_3v256x8m81  power_route_01_c_3v256x8m81_3
timestamp 1763766357
transform -1 0 25016 0 1 43285
box 349 1275 1049 1701
use power_route_01_c_3v256x8m81  power_route_01_c_3v256x8m81_4
timestamp 1763766357
transform -1 0 23866 0 1 43285
box 349 1275 1049 1701
use power_route_01_c_3v256x8m81  power_route_01_c_3v256x8m81_5
timestamp 1763766357
transform -1 0 21690 0 1 43285
box 349 1275 1049 1701
use power_route_01_c_3v256x8m81  power_route_01_c_3v256x8m81_6
timestamp 1763766357
transform -1 0 20713 0 1 43285
box 349 1275 1049 1701
use power_route_01_c_3v256x8m81  power_route_01_c_3v256x8m81_7
timestamp 1763766357
transform -1 0 42153 0 1 43285
box 349 1275 1049 1701
use power_route_01_c_3v256x8m81  power_route_01_c_3v256x8m81_8
timestamp 1763766357
transform -1 0 36525 0 1 43285
box 349 1275 1049 1701
use power_route_01_c_3v256x8m81  power_route_01_c_3v256x8m81_9
timestamp 1763766357
transform -1 0 31798 0 1 43285
box 349 1275 1049 1701
use power_route_01_c_3v256x8m81  power_route_01_c_3v256x8m81_10
timestamp 1763766357
transform -1 0 40392 0 1 43285
box 349 1275 1049 1701
use power_route_01_c_3v256x8m81  power_route_01_c_3v256x8m81_11
timestamp 1763766357
transform -1 0 30900 0 1 43285
box 349 1275 1049 1701
use power_route_3v256x8m81  power_route_3v256x8m81_0
timestamp 1764697706
transform 1 0 -1344 0 1 -3349
box 1345 3542 61604 48334
use rcol4_256_3v256x8m81  rcol4_256_3v256x8m81_0
timestamp 1765899468
transform 1 0 42157 0 1 1608
box -1076 -478 17384 41918
use xdec64_3v256x8m81  xdec64_3v256x8m81_0
timestamp 1765833452
transform 1 0 20073 0 1 23383
box -2266 -159 21704 20197
<< labels >>
flabel metal3 s 467 20858 467 20858 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 22520 347 22520 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 23383 369 23383 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 24058 347 24058 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 25270 347 25270 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 24595 369 24595 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 25807 369 25807 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 26482 347 26482 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 27694 347 27694 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 27019 369 27019 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 28231 369 28231 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 29443 369 29443 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 30655 369 30655 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 31867 369 31867 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 33079 369 33079 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 34291 369 34291 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 35503 369 35503 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 36715 369 36715 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 28858 347 28858 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 30070 347 30070 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 31282 347 31282 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 32494 347 32494 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 33706 347 33706 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 34918 347 34918 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 36130 347 36130 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 42190 347 42190 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 40978 347 40978 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 41563 369 41563 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 39766 347 39766 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 40351 369 40351 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 347 38554 347 38554 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 39139 369 39139 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 37927 369 37927 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 375 37342 375 37342 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 345 13921 345 13921 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 60018 20858 60018 20858 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59897 43447 59897 43447 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 42235 59897 42235 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 41023 59897 41023 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 39811 59897 39811 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 38599 59897 38599 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 37387 59897 37387 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 36175 59897 36175 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 34963 59897 34963 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 33751 59897 33751 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 32539 59897 32539 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 31327 59897 31327 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 30115 59897 30115 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 28903 59897 28903 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 27691 59897 27691 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 26479 59897 26479 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 25267 59897 25267 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59897 24055 59897 24055 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59920 41580 59920 41580 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 40368 59920 40368 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 39156 59920 39156 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 37944 59920 37944 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 36732 59920 36732 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 35520 59920 35520 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 34308 59920 34308 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 33096 59920 33096 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 31884 59920 31884 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 30672 59920 30672 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 29460 59920 29460 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 28248 59920 28248 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 27036 59920 27036 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 25824 59920 25824 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 23400 59920 23400 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 24612 59920 24612 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59897 22520 59897 22520 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 347 18236 347 18236 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 438 15311 438 15311 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 273 10255 273 10255 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 356 11784 356 11784 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 351 8108 351 8108 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 357 7039 357 7039 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 387 5448 387 5448 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 351 4393 351 4393 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 385 2211 385 2211 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 356 1182 356 1182 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 349 2914 349 2914 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59898 18236 59898 18236 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59988 15311 59988 15311 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59896 14401 59896 14401 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59906 11668 59906 11668 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59824 10255 59824 10255 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59902 8105 59902 8105 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59908 6880 59908 6880 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59938 5447 59938 5447 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59902 4388 59902 4388 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59936 2201 59936 2201 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59899 2983 59899 2983 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59906 1182 59906 1182 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 25571 124 25571 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 27809 124 27809 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 30053 124 30053 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 12839 124 12839 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 6119 124 6119 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 18347 124 18347 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 7799 124 7799 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 13679 124 13679 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 844 124 844 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 22276 124 22276 124 0 FreeSans 313 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 23464 124 23464 124 0 FreeSans 313 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 24732 124 24732 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 26970 124 26970 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 29213 124 29213 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 19257 124 19257 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 1777 124 1777 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 2759 124 2759 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 4439 124 4439 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 5279 124 5279 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 3600 124 3600 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 6958 124 6958 124 0 FreeSans 313 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 11160 124 11160 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 14518 124 14518 124 0 FreeSans 313 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 21077 124 21077 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 9060 124 9060 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 10319 124 10319 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 11999 124 11999 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 20167 124 20167 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 15687 124 15687 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 16527 124 16527 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 17437 124 17437 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 41200 124 41200 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 42110 124 42110 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 39380 124 39380 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 35263 124 35263 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 57062 124 57062 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 34346 124 34346 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 38470 124 38470 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 37085 124 37085 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 31733 124 31733 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 30893 124 30893 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 40290 124 40290 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 32573 124 32573 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 36213 124 36213 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 33413 124 33413 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
rlabel metal2 s 19602 141 19602 141 4 CLK
port 11 nsew signal input
rlabel metal2 s 1380 137 1380 137 4 D[0]
port 19 nsew signal input
rlabel metal2 s 21679 141 21679 141 4 A[2]
port 7 nsew signal input
rlabel metal2 s 22862 141 22862 141 4 A[1]
port 8 nsew signal input
rlabel metal2 s 24047 141 24047 141 4 A[0]
port 9 nsew signal input
rlabel metal2 s 9970 137 9970 137 4 Q[2]
port 26 nsew signal output
rlabel metal2 s 15694 137 15694 137 4 Q[3]
port 25 nsew signal output
rlabel metal2 s 35318 116 35318 116 4 CEN
port 10 nsew signal input
rlabel metal2 s 38170 147 38170 147 4 A[5]
port 4 nsew signal input
rlabel metal2 s 37720 147 37720 147 4 A[6]
port 3 nsew signal input
rlabel metal2 s 38691 147 38691 147 4 A[4]
port 5 nsew signal input
rlabel metal2 s 16472 137 16472 137 4 WEN[3]
port 35 nsew signal input
rlabel metal2 s 16753 137 16753 137 4 D[3]
port 16 nsew signal input
rlabel metal2 s 8627 137 8627 137 4 D[1]
port 18 nsew signal input
rlabel metal2 s 9499 137 9499 137 4 D[2]
port 17 nsew signal input
rlabel metal2 s 39430 147 39430 147 4 A[3]
port 6 nsew signal input
rlabel metal2 s 8144 137 8144 137 4 Q[1]
port 27 nsew signal output
rlabel metal2 s 9223 137 9223 137 4 WEN[2]
port 36 nsew signal input
rlabel metal2 s 8908 137 8908 137 4 WEN[1]
port 37 nsew signal input
rlabel metal2 s 28508 141 28508 141 4 GWEN
port 20 nsew signal input
flabel metal3 s 59416 124 59416 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 43756 124 43756 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 42820 124 42820 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
rlabel metal2 s 43959 137 43959 137 4 Q[4]
port 24 nsew signal output
rlabel metal2 s 43360 137 43360 137 4 WEN[4]
port 34 nsew signal input
rlabel metal2 s 42877 137 42877 137 4 D[4]
port 15 nsew signal input
rlabel metal2 s 50732 137 50732 137 4 WEN[6]
port 32 nsew signal input
rlabel metal2 s 51457 137 51457 137 4 Q[6]
port 22 nsew signal output
rlabel metal2 s 50957 137 50957 137 4 D[6]
port 13 nsew signal input
rlabel metal2 s 50217 137 50217 137 4 WEN[5]
port 33 nsew signal input
rlabel metal2 s 49935 137 49935 137 4 D[5]
port 14 nsew signal input
rlabel metal2 s 49452 137 49452 137 4 Q[5]
port 23 nsew signal output
flabel metal3 s 57843 124 57843 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
rlabel metal2 s 57767 137 57767 137 4 WEN[7]
port 31 nsew signal input
rlabel metal2 s 58223 137 58223 137 4 D[7]
port 12 nsew signal input
rlabel metal2 s 57211 137 57211 137 4 Q[7]
port 21 nsew signal output
flabel metal3 s 52663 124 52663 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 56021 124 56021 124 0 FreeSans 313 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 45942 124 45942 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 46782 124 46782 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 47622 124 47622 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 51822 124 51822 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 53502 124 53502 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 54342 124 54342 124 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 55182 124 55182 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 45103 124 45103 124 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 48461 124 48461 124 0 FreeSans 313 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 49102 124 49102 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 50361 124 50361 124 0 FreeSans 313 180 0 0 VDD
port 29 nsew power bidirectional
rlabel metal2 s 2884 137 2884 137 4 Q[0]
port 28 nsew signal output
rlabel metal2 s 2085 137 2085 137 4 WEN[0]
port 38 nsew signal input
flabel metal3 s 347 43402 347 43402 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 369 42775 369 42775 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 14821 44856 14821 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 18965 44856 18965 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 369 44076 369 44076 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 21886 44856 21886 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 27399 44856 27399 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 29225 44856 29225 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 25180 44856 25180 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 31913 44856 31913 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 32783 44856 32783 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 38373 44856 38373 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 37188 44856 37188 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 13958 44856 13958 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 21001 44856 21001 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 30211 44856 30211 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 31109 44856 31109 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 39703 44856 39703 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59920 44076 59920 44076 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 52323 44856 52323 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 48543 44856 48543 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 44763 44856 44763 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 56225 44856 56225 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59430 44856 59430 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59920 42792 59920 42792 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59897 43427 59897 43427 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
rlabel metal2 s 20869 131 20869 131 4 A[7]
port 1 nsew signal input
flabel metal3 s 1383 44856 1383 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 2234 44856 2234 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 3261 44856 3261 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 4112 44856 4112 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 5291 44856 5291 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 6142 44856 6142 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 7041 44856 7041 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 7892 44856 7892 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 9199 44856 9199 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 10050 44856 10050 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 10821 44856 10821 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 11672 44856 11672 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 13107 44856 13107 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 16441 44856 16441 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 17300 44856 17300 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 18122 44856 18122 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 20025 44856 20025 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 23178 44856 23178 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 24328 44856 24328 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 26375 44856 26375 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 28428 44856 28428 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 33636 44856 33636 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 34621 44856 34621 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 35837 44856 35837 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 40673 44856 40673 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 41465 44856 41465 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 42469 44856 42469 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 43320 44856 43320 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 45616 44856 45616 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 46377 44856 46377 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 47228 44856 47228 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 49396 44856 49396 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 50285 44856 50285 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 51136 44856 51136 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 53176 44856 53176 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 54193 44856 54193 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 55044 44856 55044 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 57527 44856 57527 44856 0 FreeSans 313 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 58388 44856 58388 44856 0 FreeSans 313 0 0 0 VDD
port 29 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 60260 44986
<< end >>
