magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< error_p >>
rect -34 26 34 34
rect -34 -26 -26 26
rect -34 -34 34 -26
<< metal1 >>
rect -34 26 34 34
rect -34 -26 -26 26
rect 26 -26 34 26
rect -34 -34 34 -26
<< via1 >>
rect -26 -26 26 26
<< metal2 >>
rect -35 26 35 55
rect -35 -26 -26 26
rect 26 -26 35 26
rect -35 -56 35 -26
<< end >>
