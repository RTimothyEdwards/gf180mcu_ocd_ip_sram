magic
tech gf180mcuD
magscale 1 10
timestamp 1763476864
<< metal1 >>
rect -119 94 119 123
rect -119 -94 -92 94
rect 92 -94 119 94
rect -119 -123 119 -94
<< via1 >>
rect -92 -94 92 94
<< metal2 >>
rect -119 94 119 123
rect -119 -94 -92 94
rect 92 -94 119 94
rect -119 -122 119 -94
<< end >>
