magic
tech gf180mcuD
magscale 1 10
timestamp 1763766357
<< nwell >>
rect -202 -86 362 351
<< pmos >>
rect -28 0 28 265
rect 132 0 188 265
<< pdiff >>
rect -116 252 -28 265
rect -116 13 -103 252
rect -57 13 -28 252
rect -116 0 -28 13
rect 28 252 132 265
rect 28 13 57 252
rect 103 13 132 252
rect 28 0 132 13
rect 188 252 276 265
rect 188 13 217 252
rect 263 13 276 252
rect 188 0 276 13
<< pdiffc >>
rect -103 13 -57 252
rect 57 13 103 252
rect 217 13 263 252
<< polysilicon >>
rect -28 265 28 310
rect 132 265 188 310
rect -28 -44 28 0
rect 132 -44 188 0
<< metal1 >>
rect -103 252 -57 265
rect -103 0 -57 13
rect 57 252 103 265
rect 57 0 103 13
rect 217 252 263 265
rect 217 0 263 13
<< labels >>
flabel pdiffc 80 132 80 132 0 FreeSans 186 0 0 0 D
flabel pdiffc -68 132 -68 132 0 FreeSans 186 0 0 0 S
flabel pdiffc 228 132 228 132 0 FreeSans 186 0 0 0 S
<< end >>
