magic
tech gf180mcuD
magscale 1 10
timestamp 1764525316
<< metal2 >>
rect 0 0 700 700
<< metal3 >>
rect 0 -197 700 455
use M2_M143105913020103_3v512x8m81  M2_M143105913020103_3v512x8m81_0
timestamp 1764525316
transform 1 0 350 0 1 339
box -330 -330 330 330
use M3_M243105913020104_3v512x8m81  M3_M243105913020104_3v512x8m81_0
timestamp 1764525316
transform 1 0 350 0 1 209
box -330 -200 330 200
<< end >>
