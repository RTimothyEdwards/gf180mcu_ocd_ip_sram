magic
tech gf180mcuD
magscale 1 10
timestamp 1763765945
<< metal2 >>
rect -44 28 487 46
rect -44 -28 -28 28
rect 471 -28 487 28
rect -44 -46 487 -28
<< via2 >>
rect -28 -28 471 28
<< metal3 >>
rect -44 28 487 46
rect -44 -28 -28 28
rect 471 -28 487 28
rect -44 -46 487 -28
<< end >>
